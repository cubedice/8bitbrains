��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���%��%���UQ���?6U���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍r�	�tX�)�`���$��[dm��+@ˏ^ow�Vx���_>{������6��H4ٳ�k.w�.u���ŏ|{T%�at�3������ͧdY��]]aӶ�Us�JG�DGsc2�aB�>�;�C�l���/�@O���dR�P9sid�F�q�\�0k�5k��J�|(���u����l�|���j�I�?g�f	T��i����Zߧl4���0�?�1~�x�cX`X�B%�r���7�8�.��9����/�k���hoP뫼b#Ӡe��?�F��&4%�}|x�el���7`ɝ��kN���9�ĒTC��0��`�R&.1�w��-�95�]����k?�w�>��S�@~�w��!s.��"����dLC��%��w��^m�!=�y����h�}T��nJ8�8Y�&�\�#�W��a��#�Ԗ̋�N�u���u��Uy�PD4KU7B�����<�[0YY���\�4�s���rH
>8Y�&�\�@N��B@B����n;�q�m���mi=��B�-x=�WD���4B'���S�K��i|ٓ������v9{�$W
?%x�+�� fג�� y�dH�]��/�2�-�]?�B�nI�4q�Qt!��c��<%>ì�oJ5�%,�k�W��T�٥��T�Sҥ��|E�EYZ/� c��(�U����	x]�����O���8�t��s*ո{�x�G�F�����OwꅂF�-!d6߿��b��'�� |X��M��"�D�u���lٽ�G��k�8���҆�|n���u� �(���jV%[&��\�۱��ѕ���Z�[�0�7٢z|Mߘ����g�/@�G��P�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l����2�C�b��}�@���,������0��D��L���_�L�;l��c�x�����q��F}�#��M:��;6aJVlO/�4zG&/Ӣ6����Ҽ�\�vŻ�:a��j޽����E�4.@�A ��E+���XP��ȅ&��3J��\G�Y#�u�'�'�7��r�=�����5	���]���>����C�Gظ0�����E����F��j��\w��0] b��tY��m�1�L9e.��xu	���S8��<�J�QM����2�E~9���i�d�g��U-�e�,���6+���Aݡ�Y%T��BPe.��xu	�>��l%i�-�%t̓�@��V'I�&Pi�TD��ό���.�;�~��-�fu.$�����|g�Y�'���Xw�j�7����'�\�n`��!��B�T�\ ��:E��]��8|�;�Ojz���6ޭ�@�I��w��,>����C��(R\֎u��Pm�����j��\w��0](@X~�H:0uѺ��-��(�
t�ژq���U�[��N��:�NI+���]2�y�Z鎬�����	�7 �#�#✲�@�Z����I��w��,c�A�L' �oy�
!��9b�S� 7�v�ԯ�'i�!�q�1Ig����ˉ�1�:�Ω�s8�R�	�}�����ֶ�#3��������N��;
�q�P ڨ��S���Qߵs<��7�m��+�<4��ˌ�ň��h���T�%�/ң��n�
8JA�9���$1m�dט�w��^���֮�LV����,JHn��z��p�Sg�3��ʹ�q�T�c�$�����2T�9�{uﱶ���_
�cF3�W�a,�T�~#�%�{l�7�P�H��ea�i3�|)sՀr,��>T��M��cg�P�z ��y�����,D��c2�'v�]��T�%q���h}Nw���U�m#j[5���u�L��b9����U_�+X�Ă�L�iۂj2_?.��9�{u�t|��h���\�'c_����+*�~aM�h�8���/��n(���˧�0z�cULjaGkƊ~8����\.W^�V]��}R�wX��J�W��7/đ�d;������Ga�SO/���������P}�,*�2kvQe�z�C�f�k��+ƣ�+�ه�ݮ{��c��:KY",oMG~捼�a��%"'���Xw���,D�H�p0�����dܟz>1�Pq�@��ġC���{y����x��F�U�S���QG�/dH�:2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�vsV�(�����[�ړ��D���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcd�
?ڌvWv�A��2���HF3�%t̓�@�ۅ����*���n,�d�5)��Z^ 
u�:%T2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�i'���N�����h�x�(侑�������b4�שw��@��������4���ȗ��%"%vv�J�J�3s�"��&Y��V�r���K@Nk[�r�te�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcɄ����&���IX0F�MV�ҁGG%4vkz����`���φ��<�6�C�9�*Q��7�癆cgQw�c4~Nr_�mS8<�n)�{6�U���(R\֎u�{��b�b�*%��v�ڹ߆�p�h��d��JXl'�T��~��?u��C@�|#HK��
*kB��`x��1�, �y�`��vN;��Cٯu)����bX�m�jS����X� 2����|*�`>&S�XQ�u�j�fKç<<��lp��N�DNlvr5�Dѯ���,:&�fh��[�? h�q��j��ݚ�Н��(R\֎u�{��b�b�*n��뾦�՝� s�#���k$ (@X~�H:����dܟz����{���}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ�*�6���D8C##C�K�&�a��Rg��?G���n,�d�0q�#���Q>�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�����;e�5,��y��IX0F�MV�ҁGG�.Mm-;�d=��¾ȼ\���F�`yx�>�+X�M?��y��#�-�p�݉�|�T����*qA����6\�4�@�� �-j�1tSjv������_�l)����Aɠ�T�nGHN��R���ء�I��߸��S�Ȍ�b�W<_N[h���{�`b+���Ã��Aݡ�X(�.������6soۤ$#db�i0[��-��/��?�&��J.u�$�&�V(*�O�q�p���u^�!�`�(i3��w�`L�wÝ��O�~�@}?�ggÊJo���j9��|���G��Hb� h�ҩ�jCH�d*��=����h�(-���[���}Dq�f���Ě���ž_�F�!�9t>X��u-sk,9��n�7�Y���_j����[�SRC����P�Jb�Jo���j9��|���G��Hb� h�ҩ��H����yP��C��?�T'����M?��y�!�`�(i3���ܚ��@��f�\%���M,�ݚ�Н���w�w:�!�`�(i3���ܚ��@��f�\%����(�̚�ݚ�Н�$f��_Ub�F�S�1 ��̢k���ܲ�ۗ�DCKͽ<\��1tSjv�����l��	ͰZ����XW�G�<a��o���H�RtV�^CH$�I��*�M/*�3҃�q�}���}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t`���*1(*�O�q<��?�y9�ݚ�Н�����-J2�բU�?j���4(;�jmT�#ܲ�ۗ�DC�5��t�1tSjv�����l��	ͰZ����XW�G�<a��o���H�RtV�^CH$�I��*�M/*�3�3CE'�ֶ��C�Y�\��Ra])n#���r����CH$�I��*�M/*�3�3CE'�ֶ�����B�fĉ>99��A0ok�Ra])n#��_	�������%�������&G!�`�(i3��B/�)����bX"��ͼ��1tSjv�!�`�(i3����-J2�բU�?�2h���!�`�(i3�����!�`�(i3jCH�d*��=����h�qB��S)��}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t`���*1(*�O�qԿ#��i�ݚ�Н�����-J2�բU�?���~t�;�jmT�#ܲ�ۗ�DC�5��t�1tSjv����y��lDx�_�?���&���Հ�ˤ��Pw-�h���[~,��l�:\�8��u�k#�X�I��r�$~��SgN�D��泵��Z.qO�q���f�e���M��IZz��i�ce$�q훬�LצXS�\=g(�%�H�a������~�����f_�������B�Ra])n#��_	�������%�������&G!�`�(i3��B/�)����bX"��ͼ��1tSjv�!�`�(i3����-J2�բU�?j���4(!�`�(i3�����!�`�(i3jCH�d*��=����h�'i`.���}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t`���*1(*�O�qe��0�U���>e�FW�DVx>74/���1�L�3��mJ�0�6�����1��ݘ����$�)�vx�-���΁�kk�d9�������!��<�`�s��|�;�Ojz�!��_�*9 �M�{�|L��+#@�Rh׎�no��qF%���!j������7�u?N� ;fh��[�? 'i��Ub����r����!�`�(i3���D4FFIc�	a�[2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��ߎ�	�>p����̢�/{�P�1|�o�u�/�Y����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����Ι���pG`���IX0F�MV�ҁGG%4vkz����`���φ��<�6���wFB�b�7�癆cgQw�c4~Nr_�mS8<�n)�{6�U��pॻ}��$�2p[_��dN�<@Iv�H�_��Q��b�z'hۉ)	66:�>��̢k���F�KD�Vr[/}>5��0jJ�_/�+�<�6�Q=��ĭ]�	īV�6�J�J����b����Zj���
��Aݡ��d��-��!��KVט$�W��7=��J���笺$gQy�f�ҫ
OԐ��X� 2�z���=�9��|���#o�]�ʄ�;4�zu%��XW�G�<b~*��s�
�I��J���1tSjv�����l��(�Mz�I�ݾ����]2�lـ۞�[9o�����k��^�1yP��C��?�T'����x��w�����"�on5��٪�e�H�RtV�^;�~��-�f����Ga� �^kM�ʏ����V?��Z���Ӳ��}Dq�f��5ߧE4��<�6�Q=Ґ80�)��瑨R���>&� �V$����l��M��/,;�.��1�](g���М��^������i���}	Vӯ)������7�8�fk!�`�(i3pॻ}��.�0�J�
3��Ϡeo��+�T[nfĉ>99��A0ok�����F��O�\E�W��4b����A��L��,�)n�r�(K��#)��,�c�|m��6�3�i�6��O���-&�C�U��)���Y;e�iK!���d.���+�^n=\f�5>��qb�V��jn,�_qxjzӝ���I(͂/f��Z���l�^!�%���6�n��j&b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h����^���H����b��]>���5��t��}	Vӯ)ÁB���ls)l໶�,��-��G��q���f�e�x��w�����$J�L�l:�
d��n��<f���=m�n��KS\���H�RtV�^�%t̓�@���'|Fpॻ}����}Dq�f�����Mp���N�DNlvr5�Dѯ�ũ��$[��=m�n��`>�"�on���"�":� h�ҩ�(@X~�H:����Sn/X��-���K���Ǵ,���6+���Ě����E�i�m}6O�D mWN��ܐ�}�-��cR�O�z�U���#�㔂zA���'(��h��N�M��nF��kJ2 ��b;�א �k/�ݚ�Н�!�`�(i3��b+}y[=�?��3�����4Yz�� VI Z��u�#�$IX���:�I��!�}�fb�dc���ډ���jVѭ@!�`�(i3���D4FF-�Ž�
F�'��L��quA0�e]'\gWg��	�Z�kfc�?)zni�յ[+8��r$ɓǃl[�Ƶ�1tSjv�EOJ�uxm���Bf�����'�PD�����g�Z��3��a���!@�f")u��r��oв%u�K�>&S�XQ�u�j�fKç<<��lp��N�DNlvr5�Dѯ���-����;�jmT�#{U�����y��km*}90� �p/�ϸ<��J�M����!�`�(i3Q� �_tt����˦G�����"���w�w:�!�`�(i3Q� �_tt����˦G��c�r%��I��`j!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě����ڻC�i�φ��<�6�{U�����|_e=���s�Q/a��;�`����ǆ�S���Q=-C ��U�