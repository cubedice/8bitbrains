��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}"6�l�:���L|�w.j��6��H4ي��2_)��:B!�b�ؐ:�{T�{df;���a,xh'�$k�w�D1���}����ň���x�w�Y��k��ı���$��������j��t�w`ۺ����N<��;��� B]�pE���	x]̃Dj#^Da����M�$����o��I�绯�t�z����)�,�˛D��w���旴4w�1����h���������$[Z�i��%A�a��gs|�e
�9��Ax!P����9SA��R����.���Zߧl4���0�?�1~�x�c�� ���"����j�͚L�	
o�;�i�8>'f(l����x��5�O���}@��r���7Ȭ�ϏI �ol[�y���Q\�_q_�'�i���m�}�Ć�,I�@�"|��Ca2�]вk0��}9)�Myիnň��h����c$����k��[/��ԅ1Qr������i���'d���C�0�%��w�Q�r�4����8ZJ*����	��ZHz��	�zy���i�!�`�(i3!�`�(i3!�`�(i3,-)��8�g��F�蹕�ڐ6|Zk/�/�}���1�1�ҕ�/37���E�D��`X��$D@P��f-�*��IHYH��cJė/�Ҏ�|O���4d!�`�(i3!�`�(i3!�`�(i3ɬc��WNPw-�h��� ��,/�J2���ں��)��'��8�-Zy?X��/4肋�FS�0���>E�C6?6�=B���:(̜����,-:���h�;+3�&�K5A�14P8�!�`�(i3!�`�(i3�0�9&،EB���w�[T�� TY�Iݹ�ˀ:��n�7�����O��t�sȸ�"rR!�`�(i3!�`�(i3R�����Uq9�w��Yw߿���̙	,N�Eĳ-�)�.|��]|F������sȸ�"rR!�`�(i3!�`�(i3��,�0	C}!&��[ܳ�G���������{7$0~'��&\VI`,�ʺ�;[��+$�6ﳌl��t�1��꧄�c����E�zy�զ3�0�jT ���#J��;R�S�!�`�(i3!�`�(i3!�`�(i3 ?[n�:#G٪�t6�yG�?� }[�KO[2vj���B�N� ��b�FP&ׇӭ��!�`�(i3!�`�(i30R��=�El����W\0���JY���y�!��_��0�/ᜒCX��)��h��ׇӭ��!�`�(i3!�`�(i3I����CWI�R��R���w`q��&\VI`,�$��*�z,|ފ������o������$�@�8��ˮ�ڠ��N�[�K5�����z1F~�����8h�M���W� g�[�ܣ(O#�e!�`�(i3!�`�(i3!�`�(i3�y��ă/W��G���������v��_�f�z�H�}tގ:��sȸ�"rR!�`�(i3!�`�(i3���ׂo�4�)�y��L�Di������<�FxNߡ�����Fz�!�`�(i3!�`�(i3�H�"k�j�EB����
'��(�<&���@��� 3�
2��k�B�p��mAe�sȸ�"rR!�`�(i3!�`�(i3��؆�}X�6���j\�d��'��_�]�0��zO�)�C�o8�����i��1�x����NQ[��Y���x�la��jPG���7���6�!�`�(i3!�`�(i3!�`�(i3u�+��{� ?[n�:#G}��F%���B$����&\VI`,�=JK�t���Z.�\�ػ�G�E@��j�g��o��/\k�l��p!!v*!��G�$U����ߪM3��)CSa��KlgI���7�����3m@!�`�(i3!�`�(i3��+�t2�8���]���[
y�s��;g�(ñЍBN��ç�"$�3�}����Fz�!�`�(i3!�`�(i3��p�!-�8}�����'��_�]��_��05�q��e�Ƃ�];/��������Fz�!�`�(i3!�`�(i3�*"�˪T��$�} ,`&�}�؝�T���ܜ?n昼�2#:�ֵ*&E�^8��xt��:_/�~8����A�߲wb��� ��WM�P[����(,)�=!�`�(i3!�`�(i3�B�'��a�{�ç�o�����0����(R\֎u��� Sgȼ�sʫ|H�ͩ�QϿ�ey��<0!�`�(i3!�`�(i3!�`�(i3��sƲ����e:��x���ᐜ����!���C�/�y9.Y'`f�������
��H�ƈQ�H��ޝ���'QԤ�7���6�!�`�(i3!�`�(i3!�`�(i3�7>�����D/͘B�5�35�#� "�q=i�/�J�0�)�u',�G!�`�(i3!�`�(i3�2 /��u��
���ƸtU�����*��>i�!����n,��'�\�n�~��q"P�H�oe��C��c�S+d�J�Г��f�u�����!$檦!�*��Q�`��=vݖ6�F!�`�(i3!�`�(i3��7���,�K�!5�����n,��'�\�n���t�u�?9Pjp��h���~�I��J#�2o�lS��?ꆂ�5�80�[X�b\g���J��<�i��o�]�E�%X(R�6���G<�ok��u4�w��dr��l"�X[{�25�M�1�>�J8�����È���_����Г?����."���T��� ���8ZJ*�`��Ā�	���8�� �Ļ�Q�?���c�r���q�sϻƫ}�=�������d=���q"_�v���Š~r��<Y�d��Z���붋"�M~�7>�����D/͘B�ۭ؜�J��Jt:��v{t��qS�j�e����������,[$��.`.{Xan:�ke�"�q=i%ʴ�ɒ�L��C�/�y|2I��js�B ���Wʂ҅��g�������������(��K.����M
�a��A@�r$��k���:�nj������y;�j���F���+2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE���Q��f�SR�v�����������\��o�?�m݆�8m�4|/yl}Vİ�6��$�.��Ԫ^��rL�%�7��Ŀ<Ԫ^��rL��c5����L�^
��r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!M�c�0�gB�1���i�D��0�������"��g_LG4A��/���N9D<���]ȟ!�� 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������ݧu7Y�M�+|�#��Byl}Vİ�8�d��N��yl}Vİ��8m�4|/yl}Vİ�6��$�.��yl}Vİ���Q��S
�yl}Vİ�M�W9�f^�yl}Vİ�����k0e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���2O��'HY-w�Y��k��ı���$��������j��t�w`ۺ����N<��;���u��w)�S��X3�����0ӵ�첱�)�A/4)J��ѕ���<l���9���S��9���@`��#e����4�bC��\u˻���R	j�JE�����k�8���҆�|n��1���N���	9����R<j�*�Sd,�ϱ�����p���kIFg��4�����
� �AH����eǓ�q+-��_��ƼsHcy�ߥ@�΅iG��wg�k��6비<+M�^���Qk=0Q�9o=j�+xҏ�����F������r%�<���6�|��4-�Q�,�єu��w)�S-!�����p9�AE�z,}�K;Qzd��N�Ÿ?%�b8�<�#�1-@��XѪdbm�!=�y����h�}4�1[k�8a��S����q $�^�:�Sd,�ϱ���+��!I��+�4r����C��iF �,�i!���Z��g=7W&Ş(�@ N'����f�hV��{V��T��� ���	FBX :#ب�Re������p�U�;��|BNh�m ͠c�3x��%��7�t�a�Q��щĽ��1���_����c��H�w�ǩqf�w%/B ��U�gf���^���	��'�;h�$8�k�8���҆�|n��]W Z;��TB�2��;��zoAoJ�Й�m��/K5r��!����%������&Wf�W���\�4�s�q�=Q��xjh�6g��̲��I�6�O��;�I�Sd,�ϱ�Q�%q�uS4My$y��UFt�?K��W�u�A��xY/Ų�	��
n�'���tj&J�p�J/�~8������r�O��C��0��l�3d�\`)��I���	���I[��@}c!�zg�Z�$e0���0�)�W
:�D���]�o�Q��.��&*����"E&��� ��������F�6*g^hI�χӌ������C|
r�O��C��0�����}�
��I��d�;N�%�rJ�QY!�zg�Z�$e0���0�)�W
:�D���]�o�Q��.��&*����"E&��� ��������F�6*g^hI�χӌ������C|
r�O��C��0��0RC��L���I�0�3uE#�.+;ƘP�7C��H�?*�D���;MV���L��3��eu�����F[5}%G"���	����"��y�o�+4ݒ�k�8���҆�|n���:�o�E���j:���ze��	`���ѕ������_Jp�A��)܅��r�O��C��0���df���{���哿���Fq���w�>��S���Fl��C�ըM�6�7`0еn.g��|;Pzϴ��Pez�f�{g�s�"U	�����\�4�sW c`k��TT	q��$�1	�:����Q|��Ƌu�5Q�o�F`A��PtF�.B�
m�ݕ����^z���e���C��B�"��@!�
� �AH���g���	� �b5z���lR����O<��j�4���QE���Ý�M���AQ �����Jw�)��e�0
A���l6��n�'F�H�(�/�r8@��Ƥ2���_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc$��+�{c"G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s���ħƿ�9c:��{~v_z�m%̼�ħƿ�9c�1��8�hs�R�T�ܷ��WL�C;UU����w���C3�k�����ΈIn'�J�gs�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S�7���I䟹�%H�$2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U�����ˉ�1�:�Ω�s8�R�	�}����pn�R��}"6�l�:���uq9����e hI�ˋ��vE-,b����Ǘ�Y!�`�(i3x�]�V��ι��QG���/�}���1�1�ҕ ���3�ҺIÙ=�HF���m¡Cd�_���+��;"�g�E����F�'n�^0o���˟y��)��'��8�-Zy?X�!�`�(i3JHn��z�/ue:�<� �vBX�y�`4Zp��/�����Q�^�y�zL͊�q���Vǃ���*L�E�w�̙	,N�����JHn��z�w٩L7��HUv�׿e_=����Y.�J�4�e�(�4q���ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3����j������)���g�{V�b!��u�$M�Q���?���\z-����o���������i�A( ����_ֲ��mŹ�[�g�DPp��&\VI`,�=JK�t0�`v!�����h��*��{m��=��9౲��+�J�������V����(��ؽ7$�	�s}��[	L'J����Rb��Y�W,�KYeu�BY{Y����H���/���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3i�/�
���)�����`�-�q�/��s'�\P�����i�X!�!D��(J�fŌ��P��\�v���GAџV������!���C�/�yT��H����7�ܥ��2��t��m0����r'��˝Sz��E�4.@��n̈́�zL͊�q���1m��d+0�l�R<�q��f�}��h�'f R�E����F��j��\w��0]��0�&�ͭ�h�O�0c��Et��q���U�C#/<���q�VP��@�����ɧ�J�8�J��	��	Mk�rN�By3��<�]�!����M[��Ǣ��aX� �䓒��x�O�,�j����0��G�4?�@IE�U��>��l%i�-�%t̓�@���I��gs7��-��%Mό���.Ӂ��̰�!u`Ʒ%k�����
L'���Xw��E�d��7#1=��*Yl���#�]�!����M[��Ǣ�7�]X]��@��$�K@IE�U����S8���IO,�?9Pjp��}%����͋�7>�����ǚr��y���Δ��p�T�\ ��֕ߝԀ�ح8Y��fU�aB���$�O��1���H���;��"B��$I��w��,c�A�L'Qī�*pY��am��	t���o����s����|#9��Ė�{�!�`�(i3��(�
t�������2%=dϖ�i�q㧵�0������0��D��L���_�L�3��0I}.�ANMs)�C\�?�h�	 h���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VciN�p׏.� Oag���:tӫ�C+��T���jB�Fg�Y씤`��p]�=�_ZQ�a*� k��=�R$��W��O�דW3�+��m\���X�q�E����F�_���˸@����gG��p����+�&�
�b9����`�Z�kU �o�:��7�n�s5� ���3�Һ��7U��sb!��u�}���yb��$��R�lD�]�!��	Ǹ�y85�B���0�1���U���&\VI`,'������݃�Q[R�75�e`��9|�;�Ojz�ǐ
��4�%Z鎬������_�,�[/�cWM��`�������Q]� _ό���.�}�
�?��(R\֎u����}����d�٣���N N�S�+w�7�
�p�	%6зq8�Ј'���Xw���,D�l�.E#������}��n`5�fK�\w��0]����ըi:�HCaIMl��*�>^&9@^7&ģM�I,�D�y:#9�]�B���' ��Cҷ��ecx�S�����S8���IO,���������9b�S� 7�v�ԯ��Q[R�7����n9�O�M:R	詆�����f:�HCaIMl�*;L����b!��u፪8�ܩ�ò3{NĢ:Ţ�q���U�`V�-(�qE��6I&���#���i5�S�%t̓�@��+�#i�����n,�dT�4��i��$>�c�^���!�:�NI+����	h��4��+��\��!�)HnvKr�3�͉����0��G"��������0��Gu�����ei��$>�c�kX@j�N�{u!��}�5��ę��S��!���j��A�7�]X]����,�\� ��%�D�v�l�Ū�TD����>�֔،��t�h��W+��W��7�]X]�}�4��d��D24N<I8����\.W^�V]��}���_j�Nh�EC��Q^�MY:�́# (�套�qD0Sh�Qc��/z*x�n;��|B[�x��ޗg�%���۞~��3R7�j�8`�z.1�1�N���PϾU4T k���%f/MR�V��6h���v�䩲$��<k�e٪�n��NG	�L,�N�C9*�¢�"�,�>E���,�PK����Iihs[g��DW��ԅ1Qr��[��l_ ��b�FP&s��K���!�`�(i3�i3<�f�D.`�Z���N}�m��{W`�v�L�ȱ4b��(�зq8�Ј'���Xw�j�7���7>�����ǚr��y�_��wBW��8���/���+x�r�}�9�P:��&sq�?��I!�`�(i3���7���~ֱ�q��>�L��p�T*��X�
!�`�(i3jݭ�F���%,�������;���EWr���z�щ��X�V�~h���D	��U{S��N��Tx�*aE�ֱ�q���z�␥%�"�Z1��2�A�dvзq8�ЈZ@�6������Uh1�yO�E���%�;���EWr�P�SYG�_!�`�(i3����$OV����(Q�������~�26��\��v����C9*�¢���d�������|��1�KB|1<\�~�26��\�C�LsM~��C9*�¢���d�������|��]��B����~�26��\�H,�pz�oo�@L=:�e�v4�"���Mf�{�&�t.�}��n4s1��7�癆cgR������������ h�ҩε�Ŷ�O�N��}����(/g�	�dZ#'��� h�ҩ��SSB�����B �����)P<�ܓ�Y�/��@��,�[��$�w<���x�����[	J��;��}Dq�f�3���Z[�{�]��~9��c�	?�N�����y��j��k
�X�nZ�l^@ !M��,%�R�HƁO�KLd!�`�(i3}�<?�� �o�<��p>6fs��_+L�H�RtV�^�wbk�$����$��ӝ�9��,@=ؠ�9�!�`�(i3� ͷ�	����R�����~�����$PW~.!�`�(i3�]��/ݐ�?��<*��X�
�:5A��p���N�p��8얄�Y�l,�(��vЉRa])n#���r����i`YS���{rB
�h�|���Y�l,��H��Rߧ{��d4��/��@���uSuC�hok��u4�D��'$�0��g��C�/f�	��m������G\~q~Qv׀�r�?`�f��$(���&kօ`����0`.��J��X, ؖz��'�^�����ݚ�Н��r'Z1p8u̀A�p����"�C���q(��؛�4i0��m��H���'��v�|��{ֱ@�`�7t}��p!!v*!��쬭-c�����m�����r�����n��NA���rU*��-�������}Dq�f��n��N��e9���RCJ�����ԅ1Qr��~D��!�/�o�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWNq�\E��0�'�Kխ�n��>�my$�N��{_8�Y��=�}�Vݨ�:5A��p�(R\֎u�eK�	�$V�%��v��4���kcg4�Y�J��I����~u/��kOT*qA����6\�4�@�� �-j�1tSjv��
�t��T&��ۥ`�M?��y�!�`�(i3�]}+��+[c�y��6�$��^)B��-ײ����o�N�㐜��xQ�1tSjv�X�o|36A�P%���y�TV~r�U>��O.�a8r_�=���}Dq�f��Zj���
�7ص��s�k��vy�e�9���L"�j_DK���<`*�+�lY�I���3��gCu(o?C9��\��E�H�RtV�^;�jmT�#-���H�� �5)��Z^�d��-��!��KVט$�W��7=�eu�j�~�e������5)��Z^����xQ�1tSjv�!�`�(i3<���K<�Vq�|`kK��I����<����1tSjv�!�`�(i3�SENan&���ߊ�ֲ���ܜ?n昼�2#:�^�V]��}>�C�;�����:=!�`�(i3.��J���&_��=]�RCJ�����@�ĵm�ݚ�Н�!�`�(i3��)�hV�|��L���ʭB�?�`u��r��!�`�(i3!�`�(i3=aUh������zbG�ZVٲ���<���!�`�(i3y-�S��E��*��Sx֐�M�4m�ˈk��Z��ݚ�Н�!�`�(i3?V��j�c1����?���L)��{TN��U���'��L�xt!�`�(i3�Ra])n#���r����!�`�(i3�wbk�$����$��s��K����:5A��p!�`�(i3?V��j�c1����?��&tS�D�'���Xw�j�7��Z�qҪc��(jy9d$���?�y�B���0�&�����ݚ�Н�!�`�(i3$f��_Ub�F�S�1 �!�`�(i3�� л�YJR��~6?�g �
�9Mma+!~�\R�ƨ�	a����X5b��u�0:#���"!�`�(i3!�`�(i3�HfCf�&�A��h����x&�K���q�I!�`�(i3!�`�(i3�^ ،�X, ؖz���d9=���u��r��!�`�(i3!�`�(i3���gRI/J�a$�Y JP�l��"\�$���!�`�(i3!�`�(i3��Ě�����}Dq�f�!�`�(i3�u��A�0�Ή*��a��2S����R!�`�(i31���~!�`�(i3.��J���&_��=]�RCJ�����@�ĵm�ݚ�Н�!�`�(i3�i7N�_�wDo�h�'�t�Z�f�t���p,�7�g��U-�egt�n���!�`�(i3!�`�(i3�	�vjGB�D�|�d��)��U�UH�RtV�^!�`�(i3<�6�Q=�We�
s�E�ڭ�O�q3Ȍ6�!�`�(i3!�`�(i3��O��9���:p~	E�<l���m�t>b8!�`�(i3!�`�(i3EOJ�uxm�PQ%cp��gR;#H��q�M�����ݚ�Н�!�`�(i3��w�w:�!�`�(i3!�`�(i3T�8o��7�Wp��9B���@�ĵm�ݚ�Н�!�`�(i3EOJ�uxm�PQ%cp��g��51�X�c�rs�i�}�O��LTSG��ʎh
��������n,��'�\�n)���	6�!�`�(i3!�`�(i3���F��O��ݚ�Н�!�`�(i3���"sS<���J�4�KXh��`��1tSjv�!�`�(i3!�`�(i3���Y�l,΁�a�n��]���]���1���ݚ�Н�!�`�(i3$f��_Ub�F�S�1 �!�`�(i3�u��A�0�Ή*��a��2S����R!�`�(i3�5ߧE4��!�`�(i3��l�^!",oMG~�@�S?�PmƊ��NM���!�`�(i3���F��O��ݚ�Н���w�w:�!�`�(i3;�E���Ν�}cP%��HU#;��Qz �k�w��ݚ�Н��H����yP��C��?�T'�����|�x@|�;�Ojz�$�AՁ_�mS8<�n�ݚ�Н���+�t2�|�;�Ojz�!��_�*9 �"��ӌ�r!�`�(i3q�\E��0�'�Kխ�?��ِ��E2�DZ��O`�� \)
�:qEp'{w#/ B!�`�(i3�%t̓�@��5)��Z^�q9+t�}�ݚ�Н��wӨj]h�O�M:R	���hIf��{_8�Y��M��)=໺(ӈ���]!MuV�	!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�t�	��x��ݚ�Н�0��l!������� �'���r�����Zj���
yP��C��?�T'����x��w����|�;�Ojz�$�AՁf���fa������0��G���_��8k��.ͥ�H�RtV�^4���kcg4�Y�J��I����~u���NM���!�`�(i3�(R\֎u�eK�	�$V�%��v��!�`�(i3q�\E��0�'�Kխ�n��>�my$�N��{_8�Y��=�}�Vݨ�:5A��pfĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹����:EM����Lg��h\K�5~�ܷ�S�<A"E&��� ���������^�޾F[j"]��	.�
�ɺquA0�e]'\gWg��	�Z�kfcj��r���iI9�o«IX0F�M��V8zA�|Q���м���qD��=a�^7�1tSjv�Sh�%Ͳ\rK�Z�u�Q���'�PD�����g�Z��3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l��	ͰZ����5)��Z^�d��-��!��KVט$�W��7=G��Hb� h�ҩ��H������V8zA�o��<���� ��V��G��<��
�-�ྜྷ��H�RtV�^���1� �.�
�ɺK� |�>�!�`�(i3��jVѭ@!�`�(i3��z��A�����**,n��V8zA��I��`j!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ�0��g�~�!������wP-�H1��֕q1�r�5�Y�w���
��v#�	l��lB�rq!�t�=��S[W���m�Ǝg�u-��llI"o@E �Xx�Dd�3l6�o8:4�I���c�90Mj�dL��q��É~�nJb�G ̵x�xx=�k���,� ��b�FP&s��K���,ԯ���gnņ��#�b��~�26��\2|Oo�{b��5c�;�K ���l�;���EWr��Ӓ�a(���!����iE4���9�@�*8��ڊ��
��������B�~�26��\;��B�lXFQ+��1%±�sR�{F;�f��X��2^"xm��`���φ��<�6�*$%M�֞�BW��\_\���F�`y������T�8k��.ͥ�H�RtV�^-��>lf+��]�p� �<�6�Q=Ø35�Ƞ��_�n���k9u�O��[
]&M��=���f.K���+,ꭒ���A�59�-H0V#
�@����}���yb��}-�k�D�5�q��e��u��r���n��Nh�^"�Y�.����nĞ�;@�1��i$n��Q=ߎ�����,�����l�)��uId#����*�����l��mMJ0z�}�5dg��nC������.x�[�Ё�2�Y!�`�(i3�S�Ĕ�Z�����:�\�R�w��j���{ֱ@�p��=�:uE@��j�g��o��:[q"�wP�A�
�����=@'ѥ���w�w:�!�`�(i3�GI�\�0�o�BH�n?a�ƙ˝i�����0`$f��_Ub�F�S�1 ����F��O�����@|����^a�nu4Bޗ��jw�	���|#HK������ �'����u��r����#�a�Ą|�;�Ojz�$�AՁ�Va�iryP��C��?�T'����x��w���꽤�*�����:�I���Oj�\Ʊ�������=aS�H��ݚ�Н��A�Z������**,n-��>lf+��b��~$�!�`�(i3���+,ꭒ���A�59�-H0V#Wx�Ա�%��ݚ�Н���D���l$:���k)��'�i�*ڶ�UKs,���O�޿M���$�~�}�ݚ�Н����Ȋ�?ӳ4�;Ⓠ��3��%�
�T�r�5�!�`�(i3�j����D_���w�]Jq��BѲ�+���L>!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�*$%M�֞�D��G��V]��'�H{%!��K�}.���L�Y& ?[n�:#G)Vb6^��*����(ཉ���S����v�ZT�ļm����تT4^��Q0S&",f�e�� 7��{���������m����ğ��Q��]�Q�]�(۬�~"ֶ���y��,��K�I� ����'z����;���EWr�P�SYG�_������r�Sy�n�yLjn�=m�"�2N��n�[�hŽ>톛z~$���{��m��֧�ǌo�9�(j�R$��;���EWr��Ĕō�����<�u��s$y���4�G�0�N}�m��{u��T�ߵ�sg�vRBJHn��z�3���<��;���EWr}���yb����*U���N��B�)Yd�G}%����3f��gmJ/�����^a�nu4Bޗ��jw�	���|#HK���JK���q�N�ǽ��܌��!��A/��M�Ի\1^O�LԌ|S�Fe�<<��lp",oMG~�>y�pA��x��w�����$J�L�l:�
d��*1Q\ �ޙp��ī��u�h1�������",oMG~�>y�pA��"xT��z�T/Pr
�ҙ_dW����,|ފ������o�����kL�@!�`�(i3��L���fƲ��>e<�6�Q=p�m~|�ְ��$��w��~z����!�`�(i3�����i�m����pe�'���Xw�j�7�����P�|TF<�'a��T��&\VI`,zF��^�=�*�$���i5{��s!�`�(i3t�td���5�ݓ�W�����i�2��&U�)j�S!�`�(i3kk>C�������\m��O��*�*!�`�(i3O���8z����( k��o�{��Ļ�*�@;��-b�uE9�+��!�`�(i3�P�SYG�_W-�������������>�uo"�����h1��'�t�!�`�(i3��_Ѭ�Q����%%�x�����y�7�4��}��)p��S�0�9&،��F�z�8#�\aьIR=�THIBY��v����?;���!�`�(i3U����ޚ�W�o]��e��'[+qg֚�v��?+r
K52��}Dq�f�<�6�Q=��^eY1�0S&",f�e����_n�����������"}����e����#�sDCq֌B����k$ ���y��lDM>�63��Mr�J�M�"�scX{�X!,;�jmT�#��N�T?w��l��N2B���o���%�ɍ��=!�`�(i3H�����?�@,��V�~�C0�C�(�ߜ1���}Dq�f����%>�rGO�D mWN!�`�(i3��m�5h1�^��,Q��4�7�K�ŠX, ؖz���'����u��r��!�`�(i37�:t�?S/a���X��J%�A��m}wd]]��$��'�l!�`�(i3�a�}�$�ϔjZK��#��_�?�tT�_�X�p�c�ݚ�Н��/��@��R��E���4T�Sq��{�X�p�c�ݚ�Н�����l��/f#�]h(|A�+�پu��r��!�`�(i3i`YS�������|��CK��!�`�(i3����l���J|��ȧ��lW��I�x �2a_��v��ONH!�`�(i3!�`�(i3:��kp�.,6�;�|iM�s�Ӟ*��&\VI`,9��9dJ�!�`�(i3!�`�(i3�GI�\�0�c��v�}���yb���tm���ro!�`�(i3
�:qEp�;�P�t�5!�`�(i3
�:qEp�;�P�t�5!�`�(i3fĉ>99��A0ok��!�`�(i3�GI�\�0�QWW�Z鎬�������(���Y�&�-��Oj�\Ʊ؀�o�P�}���yb���}��0�X��v�9��!�`�(i3��ۢ .���dg��z�|��Ǎ���&e`_����%~��#�8�C�	�����!�`�(i3Z��JP�����>�Q��!���c�A�L'W»��`�{͘6��q����F�z�8#3�N���[��}A?���`ޘr��!�`�(i3�: -Cx䪼#�H�r���T�:�>���g�i=:�f��&��
�>6�����YF�"�؃l��J���֨�{�Y�!�`�(i3�	��x��ݚ�Н���6���(��<7��;�x=#��la�|3k�N#_y'�H���%��!�`�(i3�GI�\�0��!���ݨ.�ϟ�7t���	t�(��<7�.���e��!�`�(i3Z��JP����wؚ���d7���͔�rs�i�}�O��L��_
�u��U.+"b4!�g��K�,>0���0��Jn��ݚ�Н��/��@��k=�E�ɟ_�ܾ7�'�� ����B��M?��=�]�֭G2�N�s���4q�.-�gg$%o�P��(
�T�r�5�!�`�(i3���F��O�VA�ڦ�c4<�6�Q=�����A��3��Y$����y��lD�鍓{�T�EB���]�(��K���'˱	��!�`�(i3� ��F�	kwJ�Rmv&&�6,d0fĉ>99��|��3�fĉ>99��A0ok��t�td���5�5ߧE4��t����M~$�)�vx�)��3�7pNf��#zP����)W�_��4zV��n|s�)>��$��|��R�3ԭ)&l�d�cG�P�U���l?��z*y�:�ly=�$T�_��2�B�1�sZ���R�ECi�dN3���Jm�W\�`!�eN#~8"�Z�Tm,��݉4G�n�?�R�O�n�6���H�V�n8�A�A�I��'��z��0���,������'n�^0o���0�yˡ�֚��IVF�\�e�}�(+;���%��e׭��,�\z�����ըi�bƑ�� τ�d�:�C/��9�PL����1$�G�͜�M�7^����1$�G��J����+��2^M���Y���wY�$��C|���NJ�K����C|�����۱������8-|�DÆ�7�U|�3�>���U��)��Ԑ#��go`iI9�o«IX0F�My�mH�6�,��XQ�$�[6{�!��6O�� "�x�H����|e"��t��k`QWf>���S[W���m�Ǝg��\+�K��~��!�������QS9>V	�����������$��N�c�0\� ��+���Y�l,V�YQ��t��t��0ã�>) c8�-Zy?X�f퀔����,>T �Jv�X�kѪ2"�ܶiv�L��k`�7�.�kU�%Rd���[�E�aV_���#�e����@ ļ�'#�э���ol#�e���ȥ��8��Y%x�&j�$�q��Cz�����WBe�R��ԓbW��)�E3	�].'�?��O�7�g�ق�𱍞3ƥB��K��3&n��T#�yY2�̾��8~e�o1n�zF(]^�Ia���X��J��W�-�`+PUy �//�����R(�4F�M7�ũhB�[��1��ޜ�%�'ȓM�Me��H��J�a�ܷ�7N	((Sb?[�Q���W���5�z5V	�qg$�[6{�!��R����D.�
�ɺ%�K��^/p�O�޿M����eo>���7]O]�|�;�Ojz�$�AՁ�Va�iryP��C��?�T'���̊�_�M86\�4�@ �i5�DiVA�ڦ�c4�I�-�}[rI:L2��J���v��tl�:�K*��gB���9XqϮ�+�N�Z�k^�U�Q��$�f�Ç{˙+�B-�D(���27:����Kf��w�n9�gg�;�?[��t",oMG~�>y�pA��x��w�����$J�L�l:�
d��o�������3��a���� 3bH2ȓM�Me��G)�X���~w�ݪ��Uʮ�V(Y%C����tl�:�K*��gB����œ��z�K�57� �N�Z�k^�U�Q��$�f�Ç{˙+�B-�D(���27:����Kf��w�n9�gg�;�?[��t",oMG~�>y�pA��x��w�����$J�L�l:�
d��o�������3��a���� 3bH2ȓM�Me��G)�X�����@p$�Uʮ�V(Y%C����tl�:�K*��gB����œ��z�K�57� �N�Z�k^�U�Q��$�f�Ç{˙+�B-�D(���27:����Kf��w�n9�gg�;�?[��t",oMG~�>y�pA��x��w�����$J�L�l:�
d��o�������3��a���� 3bH2HN��R���IX0F�My�mH�6�lZ���+�$��O$E)���t�T���S��p~����H6���a��������n@;���S&O.C�U��B��-��,1����M���K�(R\֎u����>^17Ӿ�b+}y[���̰�!`������q9+t�}��=����t��#3H�˘���o%��Y���G�&ց�*欈2��@x�3��Y$�k���&��.�
�ɺ%�K��^/p�O�޿M����eo>��J�M����!�`�(i3�%t̓�@���{z�n״$(�>g�
�:qEp:䩒=]'!�`�(i3�{�䕀��jul����l��i�	-_�����>w��-����!�`�(i3�K�&�a�W�^�|�����NM���fĉ>99��j���Gp�ݓ�W���rˬ4=І�J����+��Tٗ��
QV�H������V8zA�:�Xu��r����l�^!��'(����d�L����|e"$f��_Ub�F�S�1 �k���&��.�
�ɺ%�K��^/p�O�޿M����eo>��Hp����6O!�`�(i3�%t̓�@���{z�n״$(�>g�
�:qEp:䩒=]'!�`�(i3�h�͍��&��8�'\0�H����-� ����l��i�	-_�ވ��*I���b�Bϱ�}���yb���ؗ�l��ģVR���z����>w��-����!�`�(i3�K�&�a�W�^�|�����NM���fĉ>99��A0ok���H������V8zA�o��<���� ��V��G��<��
�-�ྜྷ��H�RtV�^���̰�!`�����'�^�����ݚ�Н����F��O�VA�ڦ�c4���'��@�my$�N��ݚ�Н��(R\֎u����>^17Ӿ�b+}y[��l�^!7#1=��*�#QSU:�����|e"t�td���5?�{�X�[�g�DPp���ܐ�}��15mo��ލ�f����`���*1Z��E��3?�d���&�i���\ݰ��x�9D�NV�h\K�5~��9}�Ƿ�J8����W�X0�,iO����qV��9`�p�0߼
�d� �!��]y�Q�'V]�<�T�bCJ�L#��K!�#n��],�W�8"M�5�O�%E#P�%t̓�@���ʳ�(�^���H> ����%�k�h�c,.J��$U	�hz!�`�(i3!�`�(i3}Y;�jn���̰�!`������h��N�M���TB$�V+�B-�D(���27:����Kf��w�n9�gg���]�e�!�`�(i3!�`�(i3}Y;�jn�.�g3Zv���� ���#qj7��p�Hs�N�*���a�*�4-���N�M�v!��$%(�jf&�~�7�;�y�>��}����e�{d����Zq��>z�����	�}���\-��U��)���Y;e�iK-pm!9�>��n4s1��7�癆cgR������������ h�ҩ΋�Q7lY��״$(�>g��̢k���F�KD�Vr[/}>5��0�B� �b���H��������0��G���_��a��o���H�RtV�^��~Щ�%��v�ډ��%>�rGO�D mWN��Ě���aT��3G�IX0F�M���]
/};����\?�u)���p�@OM.Ir���٩h�U�)3�B6#o�]�ʄ�;4�zu%��XW�G�<b~*��s�~���)��g{�d0�W� g�[��%vCчƖ��Y�l,������5���S@�b�F1Q���X��O���r����!�`�(i3x���Cr��B�%3�Y]�|�$��A
i�eL!�`�(i3���D4FF�\4�D{O8�_2��VU(��z�j�:�h�²�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ſl �