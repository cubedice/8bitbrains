��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω����	8��7���I�N<��;���Z��4d��{�
��|��Ȋ)zo1���á�K���b��j.~���m��+?��bV��ݙ���M7\F���r��C>C�݂�N$��/���	�0���'v6�o�"c����A�&�8d�v��x�۔7�D��:�b�#�Bn	����I@beB��H��>I��4�G�x4m�T
d�(b��t�켻�S���c,31�-elwB(�93;2���Zߧl4���0�?�1~�x�c,��ws�E�x��Ѭ��S���;?�jN5#��G��Qp�'���G����a�����(�I�?g�fY�~�a���+�Uz�QL�]��;�I�Qg�@zh�S҆�|n����Շ_ Q �����4��G&��GJ�Й�m��/K5r���8(�cL�.��4�����
� �AH���g���	H�Կ���>PޙQ%շ;���ӡN��v�ӫ�!NX�B�����RL�a)�ƞ��U<���H7��)5#����Nr��堅�7C��H|k�H��'js�;���"��y�s����o�k�8���҆�|n���:�o�E��c�U �=m}�R�<�3�J�Й�m�R$L=����P�X�;Qn�6
�D��t�b��M
<���٪�s����
��n�NQa"_|���voU
� �AH�)��H�]+��3�U��ڿ�e�)�fr�'�F@�4%��Y�d�u��R;+�����_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hl7�Fmi�E+���WY`�`��yZ鎬�����R�LM��ħƿ�9c�5(��}���SaB:���
�vG����BP�m��+?��bV��݊R$��������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ��,5/�c�����<��`U���/�<"��0�0�G�߲�R~�e�?��S9K��B��)]�_��mNc`A�qJ;���K����Ǖ#5�u���7�Y��]�IS��}-��j8HQ�?%{B��0B���]���~68K�}:g��ۺ�D�h�N�ta�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��(�*Lj�����'3hh��
�l>п�p=	�˳͠m�xW�g]����>/f{�� H�j�(A���"��y��J�	^�M����A��`�ˋ��7�ܥ��2�U���=9�vJHn��z�c����,XL��=d��z��_#ԠKWA�s��@
H$��jtT��kU�,�*�?X�ۦ� ~�p�o�	�a�~ۜ���B5�E̳&k	�I]����R{ A=��_�������<*�(�)TQ$|e��L��]�>
����L�]�b�֘m��+?��bV��݊R$���M/�C2�62�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcc5�e�%�ĕT�u |�f�o'
��FE��?��j��2S�u��s$y�R���� �HzX�!������s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開����� }�N��n@Kۦ� ~�p�o�	�a�~ۜ���B5�E̳&k����_/�A"�U���w�c*��o#CnH	4�3C���_����$�Qu�� ��K�ғB���	�I]���d=��¾ȼƸv��*Qx���˟yI.�	���C���&����=�g0��\����0H�&Cǣ���ZqJ*A&-�Ri�x��8<��~AN�[��-_���ݚ�Н�
ҭ�3���.��oǤ)��i�ԕ�j�R�"$H)�u�T��i�ԕ�j�����j�1ajq2�/�������� #��zG����� �#�l%��xT�q����}��Ě����E�i�m}640�RS���$
�)R�@�6�֐����o���Ȱƫw5R�z0�Op�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�@Y��g����y�4r70�-.��4���;t>
�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�߼
�d�����j�|@�� "����oH�V7�ܥ��2�U���=9�vJHn��z�c����,XL��=d��z��_#Ԡ�T��Ɓ��~�26��\�b���9�g����ҹ'-�4X�I�5hN}�m��{�a��ӷ���sf����v8��j����y��lD;�X��\�����g�X ]/����H�R�c�{2��ގ�H[i��;���EWr�'�[$t)/JHn��z��c�� N,JN}�m��{B���T�D�}�+�r1D��y����~�	�a	 ]�_���8-|�D�߸���
n�F�/���he��0�U��{Q&0�����z��Q�ye�M�8z��ɐ�$`,9�H�W�?]�U-+��H�&���_��8H�+���:=H��Alϊ��4�L�����ܗ/��@���L��PB�A��P4��tT��kU��l�m��z�KL�k|�Z}V�-��Ԣ����z��Q�ye�M�8>������`�a����t�I��cH�Z��DP7��>�������߸���
n�F�/���he��0�U��{Q&0՝� s�#���k$ �߸���
n��S��u1Z3M�w�:�50`�X���ݚ�Н�� ��Bo	�u�{q��SԖ����;b�-�2��;�P�t�5���W0�]��e|)0����n�=K ���x�?�@E�w:Ԇ���� ���y2v�W�+3_�?���cn�:������a�"�_���3���%k��)?����t}�S^ÅՍ�UsMDZ8<�V�Zs˿�}w��^z[��K�j��c���;�cT�