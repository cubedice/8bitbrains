��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��maC�S�s-\gf�N<��;���Z��4d��{�
��|��Ȋ)zo1���á-�w~��d�Ƽ(��h��mo������f���F*�#C(��$.:&R�nU���T���딣0&_���X0���2|	p��rw@	@us���)�]&��_	��u|��yq�`݊�|���"rG�
���}�\�bJ(9�{��r�H�����طǪ]������س���Ś��
��H,7���E�ջ����p��;�r�6��N����Zߧl4���0�?�1~�x�c&	��/v�߼
�d�
 O4�贅���ǖ�?xA4����*����	�f+���pB�&�zR���8��Bfg�� $n�pKJ���JI����9���j��S9�h��s��|��?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD����c���o�����0��|�hJe�A>��*�X�9���$1mt�iZ]XF���������(}y��������i�JHn��z�HKObM�^��G��^���uM�����@�b�a��1�Z���=�i��i���'n�^0o����ו���E?��`�,��C��!��pJ��H��w�1T��1��ݥU<o^.K�}�/�`��zs�]���%=dϖ�i����9�����?�Y%T��BPe.��xu	�>��l%i�-̇i�d�?�v�ј�"��Z鎬����F�71�B���N��ڧ���-��%M-�`��8�4!�`�(i3Ƣ�cP���:n##���Ψ�	�ǳ�6ϔO��)�=���O����j���0z�cUL_-��!!�5�%]���a(􆿳����^��p�n�������
L'���Xw�j�7��U����z~��6��	��k/��m#�U��_D��.V&��B֥��f���F*�#C(�š�L��]�>}|��XH��9��p#�7ڜ¸<�X����f���F*�#C(������hȧ����qcW�(u�" Oag��đ�O�v���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ږ17��_>���с�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE����#�X�HN`�K���8�8e[m��PC-��i0��d�8���
�N����wvA�qS�F_���ٱ'W�w��fD�؜�ۇ�|*����)�7 ��Ƿ��;G��ÚkW�?E-h��$^(?��"��h��w���`���φ��<�6��R!��(㽬&�p����"sS<�0�zG����ZAL�:!�`�(i3���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+{k�h�+!���?t��my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	��!�`�(i3lG%��`��ǚ��ظ
��@�U#;�jmT�#��"����G��Hb� h�ҩ�?V��j�c]���I���-%f_��m����ϏQ"j���b7�S
��n@V�� �9��1�Z���=� �o�X�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�ȌtX�IF��W���E�w�R���y�wr"�`e�R��B�.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc%�����I���%�[l��(2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���i��'{�5��9v�γ8�x���"x����O�g)�X���2�-��?�d���&���n4s1�+��uK[F�wr"�`R���;h�O��� \��W��b�[�G��ÚkW�?E-h��$^(?��"��h��w���`���φ��<�6�S�@�2�e�r&D�{E�\���F�`yx�>�+X�[�G���K!�`�(i3!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}�q�\E��08��?|�,�e��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 zM#��m����F�P�7��S��h��d\�����l����� �'����u��r���2��}��e�g��)$��K���fU����z~��6��	���`y���!�`�(i3)�{6�U��$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6�S�@�2�e��NE�]�w�R���y�wr"�`R���;h�O�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���pKJ���JI�|!�x��02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�%�8C,��Y%T��BPbvI�a�L�������	(ݖ��Mb,}!K��L힏��Z��d�G}%��Ď��J�h`���i�ͧ=ys<�+BquA0�e]'\gWg��	�Z�kfc��2���8���+�^n=\f�5>�p��9	�2�|#HK��A(�c���_G��Hb�8�u?��I!�`�(i3}�gv�oE�[��s�A>�xw'��M�v�����FK��|�H��4"?V��j�c@~~K	�dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-jېI�q�������?B��#Ɵe�*|�÷�Wе !�`�(i3L�J)���� \LÐI�q�����mJ�0�6�!�`�(i3��	�V����aٔ^?�W�<����U6�bL�QY�/�����-/a8!�`�(i3{k�h�+,�NQ��.Y�{'%sk����w�;{�'8{1�'��	�2I�R�^Ƒ���K�A�'�ݪ�򈟲�Z��*�!�`�(i3	���A�҃'�)�Բc��c��`��X�����j�5�%]���p��;�{��!�`�(i3q�\E��0KI�R�''���Xw�j�7��Z�qҪc�A� ���ݪ�򈟾�����q�ݪ�򈟲�Z��*�!�`�(i31���~!�`�(i3p�n��v{��lw	�l����;�¬pX��g��U-�e�,���6+����%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�㓔�F`#Z��/��;��|Bc����MKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�sL�:�/
e���ڝ�/&��lW"`oG&2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��P�uGA��X)5�����e�Í�x���"x����O*�������x�Y����Z��d�G}%��Ď��J�h`���i��=;L�	e�7{�.�9h����t�T��?E-h��$^(?��"��h��w���`���φ��<�6�lg�[yJ�$���Yk���'ž1�|�'����z.��W��!�`�(i3��4h�=Iz~r��V�n��dK�����fF0���2��}��D�o�&��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h�'�ɳ����Q�Y�;y��v��\���
^�ݚ�Н�:
��x�{�\��N���'�ɳ���mJ�0�6�!�`�(i3��	�V����aٔ^?�W�<����U6�bL�QY�/�����-/a8!�`�(i3{k�h�+,�NQ��.Y�{'%sk����w�;{�'8{1�'��	�2I�R�^Ƒ���K�A�'�ݪ�򈟲�Z��*�!�`�(i3	���A�҃'�)�Բc��c��`��X�����j�5�%]����ha�O�RH�RtV�^�2��}��e�g��)$�]�!��	Ǹ�y85����[��xԲ ._�U6�bL��R���~����?���=�^݊��}Dq�f��	��x��ݚ�Н�?V��j�c]���I���[�����ݪ���CyW�f�tR�wX��!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M{�.�9h�aT��3G?�d���&��fւ>�ɹ.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���\����m*>r�(�H����z��0,�턮�ݪ/�5A=�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������g�z�&���&���m��y��(<�z4G-�vN��TNm=�i�?�d���&�h}Nw���� �W/chs�]�!���3��L!�`�(i3��_Ѭ�Q�~<!��9���פ��r�3���o&�B:mn�05�2���|s�g*n{��7�4��~(��>t>�r���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ځ���$���R��9jʇ���ڮm ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcF1��_}p�MC@����<πV��_Gf���D�ݪ�򈟱i�ܰA�cTx2��R��E��φ��<�6�@a� ���N���������y�:Fa�7����os�鮊gg#��z�k�H����Qw�c4~Nr_�mS8<�n!�`�(i3���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+{k�h�+xއ5����K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(�8�u?��IlG%��`��ǚ��ظ
��@�U#;�jmT�#��"����G��Hb�8�u?��I`���*1����l��U5c��=�M?��y�!�`�(i3q�\E��0KI�R�''���Xw�j�7���W�6?���O��R�^Ƒ����"X��[��	d=�4E���b=R�^Ƒ��_uc�!�`�(i3��jVѭ@!�`�(i3D�wP�/�w��i�Wg�<πV��;�¬pX��g��U-�e�(}y��YmҐ��*V�M��nD�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6�w�Qo�Q�%aT��3G?�d���&��=���^�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc"��`V�����'/:0�쵎%��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��t�[�;����L��Vy��H��w�1T}��<+���e&nς����Z��}�
�?�bhQ����'���XwM��%�p@!�`�(i3�X����t�����\iI9�o�?�d���&�C�B*��d��}�]��K���f�(}y��2�0]�J��DB�*���NW6�6�o8:4�I���c�90�Ǘa��xB��򨙉����D�Mg�{HZ鎬����Ĺ#{��ݾ�9J�ciI9�o«IX0F�M��Dr`��|#HK��A(�c���_G��Hb�8�u?��I!�`�(i3}�gv�oE�[��s�A>�xw'��M�v�����FK��|�H��4"?V��j�c@~~K	�dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-jېI�q�������?B��#Ɵe�*|�÷�Wе !�`�(i3L�J)���� \L�1tSjv��?�Ho2�j�3�� c�)P<�ܓ�Y!�`�(i3�i7N�_ЉH�T�������ϏQ��8'嬘��lC��U*A&-�Ri!�`�(i3�ʅ���h��?<�,�-���p��U)��>����}Dq�f�HN��R���מu��� �H�0��
;�jmT�#w��ϩ���k� {�s������_�mS8<�n�ݚ�Н�?V��j�c]���I���Z鎬�������(���kO��u�-%f_��m����ϏQ"j���b7�S
��n@V�� �9��1�Z���=���VvJ!�`�(i3�����!�`�(i3{k�h�+�c������G���5�%]���a(􆿳��5���=\�gL���l���P�7� ��}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ8�vme����L���p6j�"Hs>x�'<�k�%Ǹ�!�U2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��u#a�r$	�H#4�h��@!�|w�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc;�v�-:�F|9�zk��<�r�ۧ����n|�p[Y���"���B�.G��zOEX?�d���&��@����gGY r9�=�Z鎬����$oi�~ƴ!�`�(i3V�ط�a�Lqm����ޮ��ǋ��5�ź�n`5�fK�3L��'9�� л�iS@���Ye�u�ٮ����"�� �W/chs�]�!���3��L!�`�(i3��_Ѭ�Q�~<!��9���פ��r�3���o&�B:mn��@����gG�u���k�ta�����0�]�!��	Ǹ�y85��(�C)&���lC��U�T�\ ����8w("�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л��A��ˮ����y�Cf+�����ȏ���^��p�Y��\+h|oid�G}%��Ď��J鎇~as>}�F|9�zk�&��� �WaU�?2���_II�8���8��v{��lw	���:�(�V�� �9��1�Z���=�)@����SQ��wj1���+��M�,!hޖ�A$�P������5d�`UNP�N}�m��{���q0�/)ONcx�:2QYeƈ)P<�ܓ�YO.C�U��B��-{��N�i�F|9�zk���Cw(�xjzӝ���I(͂�'�ɳ��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g!�`�(i3O�L"�
08jdN�<@Iv��nt=:��:5A��p^�ט��,AJ��w�޾�b+}y[�߆�p�h��d��JXl'�T��~��?u��C@<�6�Q=��ž�Ć�T���7X���c�}��
�t��T&��ۥ`�M?��y�!�`�(i3A�ZA��S�%]n9�hr;�H���N#!�ι�IjXT7��b+}y[!�`�(i3�R'cf���e��Rz��R�^Ƒ�Ӎ��t,��g�n�פQ?M8�f2!�`�(i3�(MXdv8��n�F0k/��s�1���� ��ݚ�Н����W0�]��e|)0����n�=�H�����qǭ%!����Ơp<���H7�I	�fb~*��s��p�k���/���q&��Ͱ0��-����!�`�(i3D�wP�/�w<eп}�����!���c�A�L'0#P�O�Z�d-�~EL%�G�b��6��	㎾��;|�5�%]���U����z~��7��:��}Dq�f��	��x��ݚ�Н�?V��j�c�/���q��/O8���<πV��;�¬pX��g��U-�e�(}y��YmҐ��*V�M��nD�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6�A.��+�W�"���V¦q��G8���e�g��)$p�n��fg�����d��R�N�a��f�b�͢�7�Kͽ<\����u��m���a{7?�U6�bL��W��_��z�ׯ�1p1�Z���=��V{C�)�߯+t9�Q��n��H�[�����l�-"�Ϳ����*��8Zn�	J���B7 Q�s֊ X���*13���'͵1���疡wgQ��@��Ԋ��,�{�����D�sZ�F��_%��VM6���ڀh�4�F��D�U��z{��̵�q3����Jm�W�u�*usp\�,�G��m.`_�j����2�NV�l�$�o��bk!�Î�]�b�y�~[�#�X�&�6��ڽ�V��(��s���𓂐Z4���bG��'��عx�J��N�o��.S$P�S�="�����:���t����M~V��	��y�3�&A��S�y�v��.�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���\d=��P@����7��\֐^�݉ 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��I^
}hI��5���e�Í�x���"x����O��GV�/�$�W�M5�O�%E#P���t�&��S���^�-�`��8�4!�`�(i3<�6�Q=y؈�&t	z���e��О=�8���*;�Kk�r}�
�?����+2-�='���XwM��%�p@!�`�(i3���#}�ΣI>]���"�L��FD���m���K*��Cd�G}%��Ď��J�?%{B��0B��<5����D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcOg ��iv��%��)�S���e�E�K�$����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �!������K���f�(}y��YmҐ��;�¬pX��c�ۛw��:0���,���G���5�%]���U����z~���D)9W �;����<rKR����a{����M���o��_�Rv�䩲$���dS@Ɵ�oB��򨙉����D�Mg�{HZ鎬����Ĺ#{��ݾ�9J�ciI9�o«IX0F�M�c�E�dE2|���PW���"sS<�0�zG����ZAL�:!�`�(i3�� л�4�>������9�@f���ʦ�/\<���tݻ�ݚ�Н�p�n���I����~uK7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(�8�u?��IlG%��`��ǚ��ظ
��@�U#;�jmT�#��"����G��Hb� h�ҩ� ��ս��	�|�O�/��kOT9�O��F�`,9�H�W�d�-���5�%]���U����z~j��AH�����:=�?�Ho2�j�3�� c��P�Q�a]v��	y'�2��7�!�`�(i3�u��A�0�Ή*��a��2S����R=q��m�3<��~�
]^�E][���-�C��7���<�O�h) �p�*���-����!�`�(i3D�wP�/�w��jJ�+�rs�i��]S���D�'�)�Բc�<πV��;�¬pX��g��U-�e�(}y��YmҐ�̓=�^݊1�m+�D8
�:qEp'{w#/ B!�`�(i3@ E���߆MC@����<πV��;�¬pX��g��U-�e�(}y��YmҐ��*V�M��nD!�`�(i3)�{6�U��fĉ>99��A0ok��fĉ>99��A0ok����Ě����E�i�m}6߸��S�Ȍ5�����/V�d��])�.�g3Z�)V��B�1rKR����a��V1�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��&2��m�e�C��J
1H�
∰����X�e����#i�CU�{C��Z<]Nٌ��c�u6t�\���(@<�d�:O���w	����h��g�H@�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�0\� ��+o#-��ik%��h�r�Bi�v�V���;AD���y��=��!�`�(i3$(��>��������	(ݖ��Mb,-�E#�����D��Mm!�`�(i3?!���l�~�y��(<�z4G-�vN��TNm=�i��
nЯ�O�!�`�(i3+Ώ1;��5�}�]���LVm��Co���ע/!�`�(i3?!���l�~�y��(<�z4G-�vN�w��;U,L��bN�1��!�`�(i3�!��pJ��H��w�1T	�|¨�l��` ���"���*�4w!�`�(i3?!���l�~�y��(<�d��������v���h�n �A!�`�(i3�!��pJ��H��w�1T����NGq���Ì!�T���=!�`�(i3�5,O�39�"<��5�{ �_�t��->��=>�Y�:pR�-�V���s�~{(��	K�+��Q�&]��_kjY%�>dc`�eE���y�C[9l%��a��31U�Y��-�E#�墙������6yT��GY�<7|'6��}������lD���7|�W�q���Ì����9���ͬ����Y�|��( $)�lj�iE�EYZ/�.�L�����