��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�����|"�L|�w.j��6��H4ي��2_)��:B!�b�ؐ:�{T�{df;���a,�|��4�Q��T�*0U1�1�:�Ω�����|"�L|�w.j��6��H4ٳ�k.w�.u���ŏ|{T%�at�3������ͧdY��]]aӶ�Us�JG�DGsc2�aB�>�;�C�l���/�@O���dR�P9sid�F�q�\��"��.,���&y�t���@N1�w�0XL�����2�U�a�6���������[m.1 T�V	�tL��	�<�A�}Q@���rah���"��yQ����D�z05��ϽE��+ST-���~���W�ZȅD�h5K��*b.[P���a�5�n��E�j������k	���#�	t�z�g�j]]�����D��ܒ[F��B����m���}Z�
d~���QK�L�$-�	BV��j`��%���˛�ӲpP�eG7ڷ�-B�"�*����	�����oŐ:J\��j�t�$*.>,xa�5��6�"
#��
�ΰg�6��}��H�F��^�'�D���3Ve���E�1�g��ȝ�0��>��R+��7���6�ړ0���Yf�4�q-H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:Qk�� h��ߖ�g��o�4��?����DNZ�j׫���?_W�\I��ఽ��`g�5��!08�tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"���`���l��r����N{a�9O��
�C�Ʌ��HW�1}Kط��4q������x��&^�B�wj$g�l�|���jWɆ&6�\]�$�n�������E?��`�,��C����-/E8�)�[���6�l�|���jWɆ&6�\]�$�n�����ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�HfCf����4�cE�D.�1o��
�p4`����J�LQ��w!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л����D��ܒ�������;;��ki!5��4��)+�[Z���M>y
��U<o^.K�}��HwL�X�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i37�_J����N��Nk%���d�Ϳ�/S����#��V$T�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3q�ɣu��ۉ�a'T���W�J'�s��4b�s��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���S�	7�i�߸B�9}.�Б����c'z=�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л��x�ҷ�������?ןuɬc��WN4�CL_܆$'<��q5�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л��dP��a�s6�Z�,��po�h0�h⤥�����	h��IB��XP���>������!�`�(i3!�`�(i3!�`�(i3!�`�(i3�po守�ud;��,4��V�;e���`���ҕH{6��!�W��!�`�(i3!�`�(i3!�`�(i3!�`�(i3Y�4Eb�������犡�&Y��V���Z:�X���<o�ĩ�U���~��	h��IB��XP���B��9i��T���K֫ �F���֦V��GedTly��鍱�� �z�k�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л�|�9I����o�u�/�ޢ��v<S�N�Ae�#�k/�z�xEQ!�`�(i3��|g�Y�'���Xw��������lԇ�-{�"�,�>E����-��%Mό���.��6[��u�V�<�nbBIY%T��BPe.��xu	�`�-9v��3�%�w�;4q�Qt!���y\���[�л���7zM#��m������5	���]���c�A�L'�����CyW�f�tR�wX��q�\E��0Ww3i�|ő����E��@IE�U����S8��y�)xʔ���6��	�\�HP@�a�~�7���� ��JL�N{a�9O��
�C�Ʌ��HW��%���E�EYZ/�矘��-n��I�?g�f&:��r-,����h��c�k�����@�&_E�EYZ/�+V��i|���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hy�C���
*P�x�v�۲=�k2Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��pq����r*+(6��l�E����F�%Z�����(	�G��^�i�<�moK��ol�� ;�ss2����p[Y���"�X��eP(�p-<Ww�I s�S����*Vx����y���;��g�2*Q=F���q/���<�7�&.��J��:����K-�7����}�쐑;�L���9��Xv7�jȯ�By�`����s�Y�{'%s�Ǹ2���;�¬pX��g��U-�e�,���6+�He�-�cI�؉P�7��':Qv?seF���+�^��BY�B�6~ [�W^b�%@�c��qe���e9 ~	R�g�,�e�+�c<c�=,����wWi:rö1M(7������C#/<���q���U�p��X
�S�9�\%��V*_�ِ�b0Q��9����ݡ�-1n �5�d7���E�Ö8�g ��L>x�R]�U��)���Y;e�iKI/B޾PԐ#��go`iI9�o«IX0F�M�\F�^��������"sS<�0�zG����ZAL�:!�`�(i3�� л�4�>������9�@f���ʦ�/\<���tݻ�ݚ�Н�����=!��9����u�Y�KG���ƒ����Ș&����Yk���-����Ί��@�=E�g�������(ӈ���m�r����fĉ>99��R�V�"�0ɉRa])n#���^a�nu4Bޗ��jw�	�����y��lD�7m�T��Ʈ+ˀa/1a@쾥~��c�'2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ݚ�Н�+�DPy�Yr� A�"W�ݚ�Н����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc6^-Yu�;�jmT�#��"����G��Hb� h�ҩ�M`�K)��v8TJ���3?���q�j\�8�E�ń!�`�(i3nD5�v�\�b�|�l<�K��u�����j��؊�9ب�ݚ�Н�M`�K)��v�^J�&t���n���"GN�^J�&t��9*�����
�:qEpCt�w#��@�ݚ�Н����F��O�VA�ڦ�c4�5ߧE4��HN��R���IX0F�M�\F�^q��_N�D�wP�/�wM"�e(&8~�$��5C�����xᐄc՘w↖V��	��y�6~ [�W^b�%@�c�xY���Ҫ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��b��T�Q5| }���А:J\��j��3�v�AQ��V��������s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�&�ȫqO8u�5ǗcV�j!�`�(i3"�,�>E���H����ȯ�By�`�2*Q=F�k�mD#V���)���6��,ڵ<�����ܺ�38��K�4V�H�%�8I�_�ju:�]i�a�*��w+J����mw_�j��ɼt���?�d���&��i۩�s���ْ5
�8�I�P�,�֘x�)�T��R�7h�����t�؆r������&Ve�!�`�(i3�l�|���j;�6	(U "#S�K�.�
.�Ūz�/>�"�Ax!�`�(i3����u��ۦ� ~�p��ݚ�Н�*�n�6��.7x4�"��!�`�(i3�:ET֤vKN��B�)Y!�`�(i3D��)����%�$A�!�`�(i3��TG���P��7U��s��6��w��'�k�f!�`�(i3"�,�>E���	h��IB��1�R�{<�!�d�<,\ͨ܉p�q��f�}���;߰�`)�΁�a�n��!�`�(i3�����E��@IE�U����S8�gY��U�v���W��_�ړ8���/���}Dq�f�\!{<�NM|!�`�(i3!�`�(i3v�ј�"��Z鎬����7.~t=� ��s�٩��!�`�(i3!�`�(i3N�By3��<�]�!����M[��Ǣ�V9_=('�����"""!�`�(i3�"B��$I��w��,c�A�L'�{&j����6��	���`y����ݚ�Н�.P̐�R
!�`�(i3!�`�(i3��|g�Y�'���Xwd�n]NْJם����"X��[�'i�!<�!�d�<HN��R��� VU+I�}R�ҁI03x���� ��!�w�#������%kRq����!�`�(i3��D��������m#p�W��	]�	�M>y
��;�?�կH��t����}�(�
4��c��^�
E�;2d�~4e$�׈PzO�e�n�^�(��.�����gRI/!�`�(i3����X=n/a�τ,�e>%����̈́�vw�aS�>
!�`�(i3����u��ۦ� ~�p��ݚ�Н��^yE⛀B��+ H!�`�(i3
�V_nu�$�F5k0B�#2\z��}�� �с�!�`�(i3"�,�>E���	h��IB��`���oX:��+��PU���!�`�(i3�E����FWA{I�Z�-"{b��~Y}J��F!��&t�ND�����l�|���j;�6	(U "#S�K�.�E�p�;+�ރ;�{��C�{�����u��ۦ� ~�p��ݚ�Н� ��ߕ!�`�(i3!�`�(i3
�V_nu�\��-��u!���ǖ�!p����nZ8����</Sn��-�¾L��!�`�(i3�E����F��j��\w��0]�B�'��a�[<�!��!�`�(i3"�,�>E����-��%Mό���.�!�`�(i3)�{� �"!�`�(i3!�`�(i3��(�
t��Y�{'%s2�ew��5�%]���a(􆿳����^��������	A�/ї:!�`�(i3Y%T��BPe.��xu	�>��l%i�-�2��}����a#�f!�`�(i3�E����F��j���0z�cUL�2�c�L��lC��U�T�\ ��&�2����wC����h�1w�0\�o�8�@If@�x�OC��q��Y}X�i��ՔJHn��z��	Dۣ��$��ص�<Ux����y�mZH֫&K������ЁK��2WIWP¸��I��'�#B��FǞ��D	��U�l>o��|�=���yp�.\��=�pe�xZ�Ư&h���}둮�z[ �}�
�?�¤Gh2�&!�`�(i3��Q]� _�rs�i��s�٭���lC��U�T�\ �͂�bv��Z�͋�V���SM0.��
�CӞD�r�u\̉�!�`�(i37s�9���o��S8��y�)xʔ���6��	���`y����X �^��!�:}Пo%�KJ�g�)}���/�#��3F����Kq��R�=xZ��j�
�iB{�Z�_����D��Z�X��kf��T�\ ��:E��]��8��Ӌ�OQ���|����Lt�2�t�d�٣��v_���Zo�{y����M�V<�'S�~�L.���P�Rg.�YP��_��Tq�'?_:[v� 5 x����y�mZH֫&t��7�M~�ۅ<����6��,�9��}�c��gCu(o?Cq��9��5�O�%E#Pd�G}%��Ď��J���i��W�o�g��GȓM�Me��e9 ~	_�nhՑP�nob���At:�)6�ȓM�Me���tk�Oȑ���Rl�Vn
*���;�E���� ��S]ȋ�I���c�90�Y��y��2�QR�e�p��ν(CmF�ln)�Xn:��N�~+�|m�N�_s�=�IX0F�MV�ҁGG�.Mm-;���6}���iI9�o«IX0F�M� ��O<�(
i�c�r�xjzӝ���I(͂�'�ɳ��!�`�(i3��4h�=Iz~r��V�n��dK�����fF0��!�`�(i3I�R7�E�g�������(ӈ���m�r����Ra])n#���^a�nu4Bޗ��jw�	���� л��E�BS�+��U�,�P!6���r�����s�Yls�<Ԍj��_�mS8<�n�ݚ�Н�,��G��z0��-���\�8�E�ń!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2�$�)�vx���za����~�&���.�g3ZE��g�Hb�.�C`S�@ys���3���L=l���ӽ~\ �r,G½��n��zfH'��!���%t�.<��X� 2!�`�(i3!�`�(i33��0���ۅ<�����B�����B:�E�hi�@��՞�gx�n�%0�&���䳚�
ca4ޮ��\4T۪��y�4�)C5�O�%E#P-�U�ڽM�T���g\��U@�!�9?�\�N���4�ۚ;e���`�ID2��E�ԇmoΖz�A\�M˩C#/<���q��&Y��V�{pў�%63��If�'¼׶�@�$Yr���t2t���k	���o�u�/-4(���H�ٗ�'Z�c��;C�f
�@"�x3���P��m@4W	�`Ҧ�׶��<�" Si^�Oґ?�&3���t��X��4tΘW���T�O.C�+��uK[Fǿ)~L�zo������g��G���*y}e����y��؎`0�H�}�	76�&�;��|B��$B����:�b��t��C����2@P��k����Q��w�п?G!�`�(i3!�`�(i3!�`�(i3!�`�(i3Ծ�|/a��po�h0�h�G��،��t�h��W+��W�{y����M�V<�'w�j���g���Q��w�п?G������[?�2�u�(��h�	r���~��n�ܫ���#Y�	��J�6Ky�QƧ�-���X4��׹!X��ǛZ;f���@7��1��+���_`��S,�{w�R���y���Aw9����Och�����ƛ���t�.�Ҝ���;��G�R�f����3a�.`Z�38yl�	�!�`�(i3!�`�(i3!�`�(i3x� ',;�J�����:���t�h��W+��W�{y����M�V<�'w�j���g���Q��w�п?G������[?�2�u�(��h�	r���~��n���;{'���Y�؂U�@p�B��p!�D�V���S����W��Y%_��̙(^���/�RvE�3HN��R��?�d���&��n5����=�r������<�L���͛2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcOg ��iv�uc�ݯ����*��� S�~�L.��� �̮��+G�މ?�[�H��bD�� t��]��hN��Ze�k�jC#/<���q��?�����9��79�4��]`*����V����&��+G�މ?�cL]�I���q�H�E� ipd�}CZv�'�ZX^�O��o�u�/��7(f	�4�"����f+>��Pk2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��Pd�G-"ұ���O�ý��i��Ք� l���E[J��:�������+�^��BY�B����葏f�f
3��^�H\�5���R�;�ఽ��`g�]C�����i�ڿ���DCEF7�R�7h�,b0V�u�Q�ݚ�Н�w�x�P���E�`JcUytԘ��dʜmT]��!�`�(i3�^yE⛀B��+ H�^,�EBj�Ւ{K4�gs��,��=�<Ί�@ŋ��5��V��(���,Wc��I�;߰�`)�@M�ĳ�@���h  �G�y
N֜�sf�?ǉ�=����>[H*k`Ë�� �R!�x�����ʄ!�`�(i3&�2����k��,�:�N�*�x�B�'��a��FD�ўB-��M��B�9{~�ݚ�Н��s�٩��!�`�(i3H��bf�?ǉ�=�V9_=('>3���T��Rz(��g�o�5�g��T!�`�(i3��gń�f �&8�,�/M�Tj!���<�ry^�=�M����FfL�[K++��d�p!c����ǖ�!}�	76�&�;��|B]}����8Sq����t'3x)'�V�G-"ұ���O�ý��i��Ք*
��10�xJ��:�������+�^��BY�B�U}'FS�j��(u�.�`��ai�2K��3�]E=����`!�`�(i3!�`�(i3v!JVʆi��8�8!s�}�	76�&�;��|BS}��X���5���
�Ƕ�W�_TR�\+�[��f	�0����k��c��gx�n�y��N��?�d���&�������y�F_���ٱ'W�w��fD�1�R��c�@N� �����˧�����b����\�'��ĭ]�	�c�@N� � ��%J%����=� ò'�����7y��<����!�_b�ȅH*�#R�J�v��6�:�bt�<�6�Q=�k;��7O�>�<6�&�c(�6k�4d�� ��9ڞ����"?��A$�P������5d�`UNP�d�G}%����3f۪�G�r��  ����l��A(�c���_G��Hb�8�u?��I���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+?V��j�c�ШT�7VE�g�������(ӈ���m�r����Ra])n#���^a�nu4Bޗ��jw�	���� л��E�BS�+��U�,�P!6���r�����s�Yls�<Ԍj��_�mS8<�n�ݚ�Н��H����&�H
�D�~z�ɕ�e^a��o���H�RtV�^!�`�(i3@ E���߂�nF���<�W�.�P�	��
�Q�}!�`�(i31���~!�`�(i3{k�h�+"���j�'fr��B�!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok��fĉ>99��A0ok��W?�;�끣�os�鮊�� ��9ڞ���zNc5�V��	��y}_�|o��g��G��ȴ.~>�@��<g$
�1d�9�r5�ۢ�2*Q=F���q/���<+��O�r!�J��:�������+�^��BY�B4��$�[��{8_��>�B���m�2��}��e�g��)$�j�=D��P�_�\AF
��|���x�>�+X����jd�	�!�`�(i3!�`�(i3�{_8�Y��=�}�Vݨ�E�i�m}66j�"Hs��^fp�/~�Cs�9`�^;�2� �S
��>ߓ�~��O�1�l��g@b���%~p�G!�`�(i3!�`�(i3!�`�(i3��mqf��x����y��E�Enk���t�h��W+��W�{y����M�V<�'w�j���g���Q��w�п?GM�ｂ g������*[wL>r~�/����ȤOa�u��KZK��\_9ͫKy�QƧ�-���X4��׹!X��ǛZ;f���@7��1��+���_`��S,�{w�R���y���Aw9����Och�����ƛ������#U|�����˧��?��'W�N��_�5�a��3�C���~�H*Qj�gj��Ν����IXt�i;�rn2�H�P�n��u�|�)ǒ�ܸ�r��%b!��u�ϓ�g�I�*B����'u��� ����.O��[�'�SҖN?�%�jwI���T%���(}���ͺ�������"���T4��$�'��h:���E����;�E���� ��S]ȋ�I���c�90���y\���$VǽO��5�~r�@&��+���_����7Pw�����&��z��`H/�φ��<�6�@a� ���N���������y�:Fa�7��mךBo�N&��+���_����7Pw\���F�`yx�>�+X�[�G���K!�`�(i3<�6�Q=��S<����K��!L��3w #�T�Z��&�2���������&��[Oթ�߁�!�`�(i3n��뾦�!�`�(i3����xSC��k���4ۏ�:��"�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")z.��W�����F�P�7��S��h��d\�����l����� �'����u��r��;�jmT�#����湡N�Ւ>��4�L4qǐ#����5{|�u��r��!�`�(i3����xSC��k���4�c�gyB��->KD��	 ���F���m¡!�`�(i3&�H
�D�h�����0� ��U�_:��}Dq�f��	��x��ݚ�Н��4���i&X��7��C�����ҧ)P<�ܓ�Y!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;��mךBo�N����5Gy���#<x����,�ǰ'�J:��XD���$�؋I~m��DL~΄gO�3f��*������j���