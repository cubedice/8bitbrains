��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����T�l䮱-�㰻��N<��;���Z��4d��{�
��|��Ȋ)zo1���á�x:��*���#�� P���ı���$����1�c/~.)��3\�R�F*}�c}��uOA�ٗ��J�$.:&R�nU���T���딣0&_���X0���2|	p��rw@	@us���)�]&��_	��u|��yq�`݊�|���"rG�
���}�\�bJ(9�{��r�H�����طǪ��v���4 #e�l(.��>��'��E����F+��T����g�"�xI+r�� 0�D�A�f�mX��1��y/P!~..�䶷	5��4�|��x:��\)�Myիnň��h����ך!�AА-suF���V�@��jy�g ��P8/�{7ht��}j"�,�>E��%�bӞk)�0�%��w��j�3��z�H8�r�(t��Vd�����%��꼸��%!�`�(i3!�`�(i3RaJ���c���R���A�0��������=6W�����<K�3�gt�6V�ݵ���������?zTz0�o��e��*�z�er���Õ������)LN���!�`�(i3!�`�(i3�?���;dW3���UWn=n�k-�;��H`��!H�@�!�[���<ilY��d�"����Gi�S�23!�`�(i3!�`�(i3U0X9�[ߒ�ڂ� ��j���r��3�N�2�M�	d�K�
����!G��o���Ѯ,>O'����4�X#�Mwn}����e�r"Dd�C�vI����:�l�5����VN�K&�edR!�`�(i3!�`�(i3��.J7h���J��V��L�k;��ޛ_�.��d)ɓ\©K�Śޫ�#��P3 9�ۗ��!�`�(i3!�`�(i3��,K0��9����'*�2��^|r u��v�<f��=WL�� _�X�m!�`�(i3!�`�(i30tYK�yPVq�|`kK��I�X�+`�^"���4���Oi5.i��A�l�	9B	�i�#fCDɈ$ɺ�������x�su~��	.��m��RVP��m?Eq�Q��fE�yӏ�E�i�dd,�ׇӭ��!�`�(i3!�`�(i3^�_�~]�=Xl|�~����m�e6؟�r�Y�}94�h�z��/��PQ�A~}��/*0�(b��g��k���M���ʜ�Jo+{)�x�=�= s!�`�(i3!�`�(i3�J܏��٢���w���,ա�	r�?�#✲�@��1��A��'gKx/அ����`��o�)Wu�!�`�(i3!�`�(i3J�Y,�~)�{lN}Q�b�o�m�����m�e6��C�/�y9.Y'`f��������L�}��xİ k�ʞ�kĶ�r:w9���י�H[��e�ׇӭ��!�`�(i3!�`�(i3����n,��>]��e��2�qj�h�7pp����2u~-��)B�Kܓ!�`�(i3!�`�(i3��&'�y����s��.���Z�!Z��`�($+����������-N��]�1�l0�)�Myիnň��h����]ߺ�`@��h�h����M����CN�u!�`�(i3!�`�(i3��7���,�K�!5�����n,��'�\�n���t�u�?9Pjp��h���~��ʍ����`���@���[K����Zw7�h[��vSZ@W�ӾQ2�Y��:�ݰ�e�M�ڙ�h�Q A 2�s��7���6�!�`�(i3!�`�(i3�e��/<9K�M>�<}ҁ�La�"h�W@	��L���:?�&lt0�ê>�ʘf��z���D!�`�(i3!�`�(i3��-���g����GBJ�tJq�Wx!�f�u�z��4�4��b�S���~��A7i�z��c�!�`�(i3!�`�(i3���7���ЍU��ń���\��p�+x⣗�C��v��g`?;W���U�W�=:	v�{�H��b/3j!�`�(i3!�`�(i3_TR�\+�[�6^Հ[�fǔ��ԆUI�S��������p����5��s�sȸ�"rR!�`�(i3
�:qEp�T���A�I�_�k�8BЧ�j-�\M!�nz��m��+�<4��ˌ�ň��h������R�뙿��M7\F���r��RL�a)2�l�f4�+��,�%���pY�� e�o�"��Ը��w�>��S9�����}����j���k�8���҆�|n����Շ_ Q +i#GBp�{_������ѕ���^�m�T��������ԉr��R�E�K����ymLj����`��j�3�����l"HP�� �Q�<�l���d��3џ1�F�Z	�����ma��}c\(�T?R,���(;�uȐ��l擛&>ث_جx�xR??���\z-ܘ�u}����!�`�(i3x�]�V��\#O���oY{Y����H��c%�ݿ�;�uȐ��l�ɘ��9�GHmە,�)	�8VK�>U#4(������������˶?��xBc?	7�f�7�~?�_�T!f��\����l�����[�ZJ*�97),J�l�/�4ќ{K�!v�0`�z�4/H�49U��љ�S�?=g���9xsjɇ%�ꤸ����O�!\�/wy$�ն���z�?%B8��2<o�J���_ r��r0l8�fQ�q�tb��JD�=����֧D�EM���
+����rϓ�g�I�*P��*�C�؞ �-:���xE��� ��P����RL�a)=�y�~ ���H7�14����ؑ(�3K8��!�zg�Z�$�̹�d.ň��h��U4T k��ko�Y��6�ʯ�R<m[�Og����n�ö�4�*x2 �Q[1I�����w'�\�Q�3M���e�t��yn�	� �x�m��n~�q({L�51��;����'��%Ճ�86���H�aF��6��I���j�r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�=W�֯�ZW���xF���慼|~09h�i�;���6�ӫ� n[)Z�Μ._^���#f�EdY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc~����������0��D��L���_�L�����J]5+a�#�$�@%�9���$1m�ea�;y� ����t��=l�)��%�0|]<w:�"�,�>E��4];ˍH�w�����޳x G����^������f�j�����=6W������E����F}�=Ll���o�����[�g�DPp������=6W����,@)=i��i�����8�TP��e��� �ρ56����RVP��mA="�����9+
�����y��[�~#��#��w������!�؟�r�ԝ0Xz�#��b9���A����
�)馢䃒�t�rZ�?ђ��P^(����gi���$R���b�>�oa.4���t$W�<	ݎ�T��ߞ�����i�зq8�ЈR���b�>���d҃!�����4X%�ٿ�����c��N�wC����<Ӿ^H��	x�]�V��\#O���o+�:#�����)N�E�3��k'�r�E����F}�=Ll���o�����[�g�DPp�˜�?�������gHucN�pS��Y}�=Ll���o�����[�g�DPp�7>�����ǚr��y�N�pS��Y�'n�^0o�ՔҬ%��؍��R��j�.(Wx*�_F�k-��E����F�ҋX����>��l%i�-��E/��F�/(A=�k�]�!����M[��ǢK�h-L���H�B���5�¬����"����N�By3��<Z鎬����A��:6])���^�Va��O�MJvx�W�D߫G_"�|�2�o��C!T*�q���U��ݯ�AJם�I��gs7<��z��}�\w��0]��-K2Y���.m��
S�)37J*u>����C�Q�rG�LNN�By3��<Z鎬����A��:6])��k�{���*��� ^�e�n�� ,7�,�䜑Ḑe�p���,�䜑t����=%�G��B�p[|C�ɜi�M�g_��e۳��ZS�)37J*uc�A�L'��~�2�?؟�r�`U���6�˝Sz��E�4.@��/�G��x�8���/�I<��fҹ�\�<�dQ	���qk�ZV"���:��#tC�|�P��Х�]��:N��;
�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h}|��XH��9��p#�7ڜ¸<�X��/~.)��3\�R�F*}�c}��uOA�ٗ��J�����h�L�;��"�r�C$�q��T樞�&�P�b?�F���ȡ��b�2T��}5��W�7�pIS2c��Un�`�n��/����֧�$���xK��D>��A.tKa�;q(�I��h9���v"c'��ɿ&0J7w� a����c4d꽇��DT��8Jp�m~|��pͧP�J}�a�\����%�֒7%�\b�Up�rP��O�6U���idf@�x�OC��b�7�xة䧞4�ڕK"�hs؏ 4�+�{_8�Y������I|��0����|�9�H�d"ֱ�q����q!�[�l�M_p��'���Xw�j�7��,�\�I��U56=����[Q����Y����I	3�ֱ�q���5��99��/���|M'���Xw�j�7����rI��V@�}ݧ2N��n���?���^�:��Y�*��P/;D���V�o�7�_��$�Qu�g��-����Q]� _�rs�i�����\�k(n'A�8���8-|�DH�%�swUp�rP��O�%2����$u��r��R�@�6�֐��T��˩������H����/ʸ��,�c�D=��dv�h2kC��-�������M$��v�@����b�z'hۉ)So�jQ�ŗ�	��x��ݚ�Н�����$K7͍��hB����G�筬���[�T�!�`�(i3��$7A�fm;�O�y=شѧ��v��HN��R��bP�63Z�t��-����V��~\��! c�A�L'[����Í�4W��C7�%M��أͽgF"?�"g�������Yk���֦?ɖ��h��x\y�<a�M�4������<&�}�V��ݚ�Н�F9��k�~H����!�`�(i3�av��%7�&~e�e��E{��h޴o'
�X���|e"ʁ���Mյ����+�	Ղ�I8�y\��S��z�p��T���!�`�(i3U /숇�m.V���Q:-�;S5b	��T�.�<̎��_��6����~A���U젩`#FW8�	��(hc�)�"��}Dq�f�G�&ց�*涑�K�v�n���}���S.�3����/�f?]!�`�(i3pı��0��[�Ez|�фZ��3��w��\�W����5���ݓ�W���M�i�s4�0 L?ஹ�%�����CCe��ݚ�Н�(*�O�q4؂C��[}�N�`2���K��޵J�uc!�`�(i3��p����&~e�e��E{��h��9Z�2�"���|e"ʁ���Mյ�A�Ɲ��	Ղ�I8�y\��S��z�z�����Qn!�`�(i3U /숇̽�2,5��-�;S5b	��T�.�):�N����6���PfL���U젩`#FW8�	��ܰ�~��؜�}Dq�f�G�&ց�*��{�![�+n���}���S.�3����忝a;�!�`�(i3pı��0�������� �Z��3��w��\�W��Hs�o²�ݓ�W���u����q�t4�0 L?ஹ�%��q��=G�j��ݚ�Н�(*�O�qng5�}�mc�[}�N�`2���K��
�Ɗ-�=�!�`�(i3��p��AZ�&����`h��E{��hS��CY#����|e"ʁ���Mյ$��Q��@	Ղ�I8�y\��S��z�B��0���!�`�(i3��4�CD5���}Dq�f�fF�5.]����}Dq�f��y�"�V����譬$f��_Ub���uQL+��߼
�d,ܕ�21��IԞɹ�}�
�?��@�/�.��B��+ H=]A��O�T�ҹ'-�=l�)��%�� 	��k��#��5MʶE ����0*@$`��)^�T�H����d�٣��v_���Zo�����]��O�M:R	�G�L3cfi����hD�v�l�Ū�TD���)T&I2WM�vT�V��|�������c�A�L'��~�2�?�B���N�gl��ܬa(􆿳���2����.��DP֞ E2�DZ���PZ��8��"�7ϫ��*�.���`�������H9��p#�7ډ:=^�=��?�g�˖���R'cf��i�X!�!D��(J�f�w]�IB[�)����]�5�O�%E#Pw�����A�#���Q�X[[kl�JFi���Y�v�����Ho��'�\�n`��!��BBaYz+�Z����~R���1��� ����P�7� aT��3G?�d���&��R�7ʌ�J1����?����^��x�=WU`wl�o�l���hLI�	u)3̩W�G��!?�d���&�05�2���lO	"�����S�Ĕ�Z�q	�R�ML�p�Nģ�Z�8��D���p/�LL�ҏ!�e186?܋܇�h�'f R�U���e���`D�����Cs�r�����/���	􈸓��-�F�\�h�b��B�i��s��t$L�����(TfSW!H�q�j�iT�s$ć.&,�*�G ��@!�D6H�
t�@����~.���gɄ�6�o8:4�I���c�90j�L�A!�@��v{�G݇���6@��a]W���\!�`�(i3 �7�Q=�y�n�:ڑ�ۍ��[�k(���V德�6-���_Q~�O}+K�)����a���}�9�P:��&sq�?��I"�,�>E���2,��T�B���]}_>��J8�c!�E����F�Z�>)��oz��KUq����a���s�*�I��g�W����Q�S�ʆ�In��t��}Dq�f� ��b�FP&P"G�wk�\����b9���1]�?���N}�m��{zh��ʊw!�`�(i3=]A��O�T8�G��oBߓ��A}:h:
���9
!�˝Sz��E�4.@�o-�!���H�g��U-�e��,H/��N}�m��{�
i�F}�W!�`�(i3L���`H�j�7���7>�����ǚr��y��CyW�f�tR�wX�՛���a���H��9'p���y�x(�E��*������m� w����tq4��}Dq�f� ��b�FP&%0Z�M��L��՜-)��±�sR�{F��JG��<.+6J!d=��¾ȼ;�jmT�#F�KD�Vr[/}>5��0�B� �b�Ъ���l��t$�:�r�@u�ÅǷ�B� �b��!�`�(i3E��\�����۪%Nk˹@��]��ñ�o
� /G^�̲Q������4��G��RV�N�'�� C-��&�X��r����Ҝ���wM%���J���2o�A�g%"��/8�Nw~���I,Z��0���f���Ն� ��%�D�v�l�Ū�TD���7��y%%9���.:��Q?M8�f2!�`�(i3�JO�'����"@wOД\��Y�� �Ξ[�s��\2��Tլ�����![ĵԝQ&ޜ�}Dq�f�HN��R��Gu�"�0�!�`�(i3{[�ב�C���#�'4v~9��c�	?�N����!�`�(i3U2y�T�2U���2��&�t.�}�ݚ�Н����F��O��ݚ�Н�t�G�����DZM�J8�c!����M׮� л��ݚ�Н�E��\���Ft�[�����:�JK�2D��MY�|<NK�6��}Dq�f�1}�ั):9��tf��!��Ϗ�2�ed4���Ȝ�}Dq�f�^ &��� t�rN)X����Ȋ�?ӳ4�;Ⓠ�X/�7�D(4'H�]����_�6O����Ȋ�?ӳ4�;Ⓠޕ;j�j�������"�
�T�r�5��� л�P�|���9��V�91}�ั):9��tf��!���i��L��G_"�|�2��v�9��a3@��[/�L��O��p��?z��t�g"m�	�uE9�+���~���U�؜J��v�W�Hl���̋mϏ��Q6~�{W!�`�(i3J�����9��tf��!��Ϗ�2�ed4���Ȝ�}Dq�f��1Ƈ��,,�3 l���6������S>�;�u��tF�{F#��� � � ���ݚ�Н�E��\���/C�Z��[��y�x(��dqܧV��ݚ�Н�|��7�u�ci���{2a3@��[/�L��O��pg��`�t�E�?:�^���v�9��a3@��[/�L��O��p��?z��t�g"m�	�uE9�+�廻��j��y-ʲ�}��6������S>�;�u��tF�{F#���'��.z��6������S>�y�-�RJ5Y�bv�N�ԑP�מ�����y��lD����g���-S�!�`�(i3�R'cf��i�X!�!D��(J�f�x��2�+�T�\ ��[��(��!�`�(i3����0�������ߺ��8�ۦ�P�X��P�������pC-��h�>
A��%�.MB^Ms\HqWU���>
A��%�������}� h�ҩΉ?�W/)G0��#��#c���܎�Aa4$�+�3�t�.K��ߎ�x��y��v�9��!�`�(i3�JO�'��a�}o8g���?�!�`�(i3t{�lPz��˝Sz��E�4.@��:u]R��GX�Z�X�W�NY���eb��D@fQ�ce�c��)=�,J�� ��C���Q�ce�c�Ԛ�-����!�`�(i3�g��2����͆���_�=[���:�HCaIMl�T��G,���ݚ�Н����Ȋ�?ӳ4�;Ⓠ�!����}�:5A��p�Ra])n#����m?�V?��?s���9qj�xm�N�e�{�W!�`�(i3|0u��\���.ޟ���T�E���U�6�'�)�Բc1����?��S(�`�ՙ!�`�(i3���F1������$��;Ε^���3$�J�5'!�`�(i3�k��^�1���[�a���mk��T9s*�s}��[��-����!�`�(i3��>��lJ)�W�=�k�Ҟ�#�>�L��n��p��b�Bϱ�:�HCaIMl�i;��B��}Dq�f�`
 ֢��؜J��v<�8��k��vL n9-�N
�T�r�5�
�:qEp�;�P�t�5!�`�(i3E��\���/C�Z��[��y�x(��dqܧV��ݚ�Н��?�JY�)�q��ڍ���F1��kټ�b�	�RCJ�����@�ĵm�;b�-�2��;�P�t�5W?�;�끂W"�P�K�׶h����z%�o�{�w�R���y>��yС`�&zk8��������0�"��G�K�I� ���F�Ҡ��q��É~�nJb�G �!�`�(i3$�xKw�6��/B����~?H�?�����3@�4�;Ύ�@�ֱ�q�����2�w�]'�-Q?9��E����F��K�J���N}�m��{�K|����}O�6�T���M��VK ���l�;���EWrr{�"���!�`�(i3jݭ�F���%,�������;���EWr~��*i!�`�(i3jݭ�F���%,�������;���EWr
Cj�R[z�����/�jݭ�F���%,�������;���EWrAԢ�a\���*e>�{JHn��z�3���<��;���EWrQ�^���!�`�(i3x�]�V���ɱʊ��7*�/�. "o�M8Ԝ�������Y�W��	z2��Ň7\x�*aE�ֱ�q��(�_���ߦ�D��.�E����F[s�9�-n���~�2�?�B�����lC��U�T�\ ��yO�E���%�;���EWro��%��jCy]vLjݭ�F�����o�m�H��+x�r�'���_�)������X~�E��*������m� M_>�nݥNGz)��.��|ȃ��d��JXl'�T��~��Uг�|<�@�O�����>[�@2Y�6�x�T'_�>[�@2Y����,1�;�jmT�#��"����G��Hb� h�ҩ�f��ZW���m�F��#o�]�ʄ�0c �)��l:�
d�x{^4��*m!�`�(i37�%M���6Y ��؟�r����ڵ�a(􆿳�Εq�8!�`�(i3�#���`���@���[K����Zs��$�Z�܌��!��!�`�(i3
�ɥMz�j֓�D�l�t�Z�f�t���p,�7��y'�Vq�|`kK��I�������pp�\ì��!�`�(i3�Y闹��5�x����VY�+��I��0��Rj/�u��r��!�`�(i31}�ั):9��tf��!����WBe��XpbJ��>[�@2Y��[�[@�B!�`�(i3a3@��[/�L��O��p���F�<g"m�	�uE9�+��!�`�(i3�5ߧE4��!�`�(i3�Zj���
�7>�����ǚr��y�%�!��U]�ߍ�2d��3џ1�F�Z	��;���P*��g��It\$�ݛ5�CN;���P*e�{�W!�`�(i3.$����0�*��D�x�=l�U�-kO��u�:�HCaIMl�i;��B��}Dq�f�!�`�(i3�JO�'��a�}o8g���?�!�`�(i3�k��^�1Jbk-����'�\�n1���R��뷅Kn�;F�Q��s,�~TM�e�w�G�U�s&��*0�uYOs�ݎ�T����U�s&����\W��N�!�`�(i3�Dd�\���؞�W�}�:�c? ��@2A^N�]|-&vY��;�!�`�(i3���F1������$�ӿ�F{ј�^�ݚ�Н��Ra])n#����m?�V?��?s���9qj�xm�N�e�{�W!�`�(i3"(<K�'PyQ���4��}�@���_rS�b�8Z��W�6?��O�M:R	�گ�����ݚ�Н���6������S>�D]h����yQ���4�uE9�+��!�`�(i3����١�$�ݛ5�CNTף�[t�����������G�R�u��r��!�`�(i3��>��lJ)�W�=�k�Ҟ�#�>�L��n��p��b�Bϱ�:�HCaIMl�i;��B��}Dq�f�!�`�(i3�JO�'���Q��\{9
Cj�R[z�!�`_q�!�`�(i3$f��_Ub�F�S�1 �����l��#�X��C����Խ�TЃ�si�ݚ�Н���6��b�8W�wo_V��U'��Cq_c�!
�T�r�5�!�`�(i3��jVѭ@!�`�(i3�Jo���jQ�kŕ��QzM#��m�<�6�Q=*qm�U��g_WԽm`�P^��ݭ%�?�p}iBy��R<�pc!�`�(i3���F1������$�ӑ���n,��>]��e��^���!�`�(i3HN��R��bP�63Z�t!�`�(i3�5ߧE4��!�`�(i3�u��A�0�Ή*��a��2S����Rq� dr�+6V��\"��C�/�y|2I��jsi��3�a/� h�ҩ���6��b�8W�wo_V��U'��Cq_c�!
�T�r�5�
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b�z��O��r��s�yk<Y�
�
���J��V�quA0�e]'\gWg��	�Z�kfcM��fZ챺�k����q�hgv�~A_x^6l8���x�;���EWrr{�"���,ԯ���gnņ��#�b��~�26��\2|Oo�{b��rA���oq��WX ��b�FP&�&5�/hеR�աuΨ�KB�c
5Xn�DIc�&5�/hy�b�G2���+�^n=\f�5>��I��|ij��"�T�\���F�`y������T�8k��.ͥ�H�RtV�^d)ɓ\©K�Śޫ�#Wx�Ա�%��ݚ�Н�m#`0ً���x R��9�U+˘n����q�hgvvC���m+w���f\P��]JP3�)x���=��:5A��p�x��8<�k�e�Y�&5�/h�͵G �T� h�ҩ�m|^�XlF �%�:���Y6{��G奄d}���5�#ϙ�s��� ���G����:[q"�wP�A�
�����=@'ѥ�$f��_Ub�F�S�1 ����F��O�����@|����^a�nu4Bޗ��jw�	���|#HK�����ӪA��1h�'��H���b=�W!�`�(i3L�J)���� \L�1tSjv�����l��]�3��$�Eʨ�`N/���US��W����E1�����u��r��!�`�(i3%ʴ�ɒ�L��C�/�y|2I��js��'Q�:�H�RtV�^!�`�(i3=aUh����I,�D�y:#9�]�B�,)g	�{  ���ѡ=��mva��!�`�(i3�SENan&���ߊ�ֲ���ܜ?n昼�2#:�^�V]��}>�C�;�����:=!�`�(i3<�#��/Me�T��2:�)���/}�׏)#uE9�+��!�`�(i3mv�%�3�]-�e��v��ʡ��
���,��;�b�0a*A&-�Ri!�`�(i3�/��@����}���rf���fU�1Q�\��^����!�`�(i3!�`�(i3fF�5.]����}Dq�f�!�`�(i3T�8o��7�Wp��9B���@�ĵm�ݚ�Н�!�`�(i3���L2r{�"����N��Ưb7�Q�^8�bL�1p/-��N�]|-�}k���!�`�(i3�/��@����	X%+7U�i�#!����P�>�����T�8��dQR�?e�F=�꤇�{�l�	z9�3OK~�hGրu�%���K����4q�.-�gg$sf�e�}s��������t����>PQ%cp��g�i*�;�wa'����\�f"������WBe�IU�A����ƧG����]�w9"xy�b�G2!�`�(i3fĉ>99��R�Q���~��p����!�`�(i3��jVѭ@!�`�(i3����Q�7}Y�Q4��6��k���ݚ�Н��/��@����}���rf���fU�1Q�\��^����!�`�(i3�ݓ�W�����o߽�..f�پ��gp4/j��ㅑl��o�����zQf!�`�(i3�/��@����}���rf���fU�1Q�\��^����!�`�(i3���%>�rG�E`���!�`�(i3f���Ն� ��%�D�v�l�Ū�TD���7��y%%9���.:��Q?M8�f2!�`�(i3�wbk�$����$��s��K����:5A��p!�`�(i3C�7�/�)hL
��C��Ͳu�d�9�(�%���]v1�_ُE2�DZ��+[��P����	X%+7U�i�#!����P�>�����T�8��dQR�?e�F=�꤇�{�l�	z9�3OK~�hGրu�%���K����4q�.-�gg$sf�e�}s��������t����>PQ%cp��g�i*�;�wa'����\�f"������WBe�IU�A����ƧG����]�w9"xy�b�G2!�`�(i3fĉ>99��R�Q���~��p����!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�I��|��8������L6�>P�2-i_m�;Y'�V!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��F