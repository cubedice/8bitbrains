��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�>���U�_�4�0S�����x$.:&R�nU���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍C95^T��6\Xa��7��Į�N��=i�@x_\q��oGo�Z�������/�)��ɖ`ۺ����N<��;��� B]�pE���	x]̃Dj#^Da����M�$����o��I�绯�t�z����)�,�˛D��w���旴4w�1����h���������$[G��m$�;�`��v��p�㈍x���t�켻�S���c,31�-elwB(�93;2���Zߧl4���0�?�1~�x�c�>j����d��S�W�>��Q�d����t�mR��:�����-��3���7�Jk�b#Ӡe��?�F��&��q�©�����<�������~s���^���h��~�a��9�ĒTC��0��t�z���� �Z��[H� �?��Y2oB;sѱE�%2�}���3$�" ����f����m�!=�y����h�}�BK9�H�N�SV [?�f��%�Y�o?�M��;]�#>fS�H��K��l��fu�Z��"R��Hv�|{")8�*I��_YLw@�H����>8��\�����^gF���0r	+2MWm�Q� ���,�Nk��6S�䥭*����	�z�}ݢ�Qy�?3�Vǡ9���<aDK�^�aum�Q� �8=��,�}����;�P���Ħq�e�����4�})����_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3ts�JFAa�ߖ�g��o�4��?����DNZ�j׫���?_W�\I��ఽ��`g�5��!08d��q�G�+��T����oGo�Z�������/�)��ɖ`ۺ����1}Kط��4q����S��Ǵ��BR�^Ƒ���E����F�Z�>)��`�U+�PA����Kp&�@���k�������5	��{�OF8<z,Ҽ&���L���g���x z�Jm]A�/����<.+6J!�t���\�W+�[Z�����+�J��U<o^.K�}��HwL�X�p��76,�/^;؊��^:#�^)w�<�_Nh0iMAͽφ�4�e��gR� �ұ!�`�(i3���D	��U�l>o��|�,+$\�M��wF4��0[����	��N�Ae�#�̲�2�!ڢ�{l�f|��rs�i�� ��*b��0��E|�,�CyW�f�tR�wX�ս��Mڷ��S��'�?�]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�eן�-�Q�Z���S�|Jc��Et�Y�{'%s��.|Z���I7��-5��6��	���`y����ꢤ�Og�ś� ����]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�eן�-�Q�Z/����o<��z��}�\w��0]Y��
�iC�o��C!T*�q���U�&��GE<�N�By3��<Z鎬����y��|�!�p�tN2s���(����5���ռ�j����)w�n��ukh��Q��ņD^�NË�����8��z{��E�EYZ/�矘��-n��I�?g�f��Qө}�8o�C���7I���ʊR$��;g��4��s;�s��&<�w�п?G��q8h�G[�� 4&Ƒ:2�c<�^<�H�U�YQN`V��	��y��2����8��`+S6E���7-K����}�)��E�d�-���geW���w>��Y��$1&ODQ3�z�sis@�����]���ϸ��#|S������3[�u8�J�a3mPy��>/' k!�`�(i3!�`�(i3�X;p`�FJ���f�?ǉ�=�����hWK{m35%7� ��yDg!�`�(i3�X;p`�V�׍A�f�?ǉ�=�����hWK{m35%,�!�H<�!�`�(i3�X;p`�V�׍A�f�?ǉ�=�����h�? "a��Q�V!�(�!�`�(i3�X;p`�V�׍A�f�?ǉ�=�����h�? "a��%}w�dN�!�`�(i3�X;p`�V�׍A�f�?ǉ�=�1_�
774\51�]2�t��MJT�!�`�(i3�X;p`�gR� �ұf�?ǉ�=�t� ��O���}���i!�`�(i3!�`�(i3�X;p`�FJ���f�?ǉ�=�$�V��bst�N���!�`�(i3!�`�(i3�X;p`���z�����2� ��=�<���� z!�`�(i3!�`�(i3!�`�(i3�sg]�_�}F�r�f�t��5Z�����N���96!�`�(i3!�`�(i3!�`�(i3���I�=|�0��E|�,���6%�az\�m���Iϕ������z_۬=�!�`�(i3�&8�,�w�Qt
����+g#>�2Y��kک��4�+/r���G�6!�`�(i3!�`�(i3p.0��I�![�Do�9�ݚ�Н��5�w�yzwz!�
�W@!�`�(i3!�`�(i3���K�7��u�mD������$��`%��nx{<qH�~�!�`�(i3!�`�(i36�ŏ ���.��?e��q�9�ͭ\�j��fxj�9�t�.܉giIE�!�`�(i3���
�#1M5����yA�y��j��k��V��e�LtW��e���d�tAAI�O����0�8Xi�fΊ�}M,�d�X�N�� 6���6���0@�pgd@!�`�(i3!�`�(i3!�`�(i3xj����R��á�~O��&�C�/#�n�%G2_�ĉ�j!�`�(i3!�`�(i3-��A�sxW�O�,��L����6���ʛ�M>#�!�`�(i3!�`�(i3!�`�(i3���u�UgF˯�+)��&�C�/#�n�%,�Xʚ@h!�`�(i3!�`�(i3-��w¹��<d�,��L����6���_G��?u:�L��!�`�(i3!�`�(i3w)����*RN�]�5'p����nZ���t��˳3[�u8���9K��r|4�:���m�
��,!\4L$ֵ���A��)}���/k߬p<Y��j3�� ��ݽX�Q�L����'T���+�n[���/С���?�T!?��vSƏw0��|3�o�%,�2��E�\�tP�;EOJ�uxm�)7*{��C���C�,�4��؟O�,�Xʚ@h�d�)bU�x1�~g_cId��V��	��y��2���,���H%�Rr�����_�4u��