��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lV�t�[;�Z��4d���Ġ���딣0&_���X0���2|	p��rw@	@us���)�]&��_	��u|��yq�`݊�|���"rG�
���}�\�bJ(9�{��r�H�����طǪvWa.�U4�,3���\.�"�K����u����l�|���j�I�?g�f�;K�y��rk�gH�I�6�"�Y!����Y�f��a�Z��Vv�c
�����R��Y���`z�X���#�ӓ]����?6zՙ}�WNg�k�-i�ʓ��	�[	r�7Ѣ��K����@�_3pp҆��V���Ї��?L���u���{������`wi����Q��Բc��7_��+��׃-����R�xTGQ 6jy�u_Ĉ���rl?�4�ʗ�C��JuG"�/��m
>Qo�n<�!+X��Q:�"��!�"�^IM�om\��(&9B:���Z,��3��Đ���xΕ���}Q�Y�:��^������t����$���ӧdR�`�����֞��� �js����vb>8��Cru-��-׎"���f��sVh�a�ei�P�?�_��,�Y��oT��_�n�q5�W�@����΄~����p�H�^�O9.]`�GMG�2�3Ӭ��;�Ӏ׬V}A^�� ��!w����qz;@̉���ߊ���7/��� xJ��V�	���
��J=+J4J9�B_q���v�p�*��	��6Ǯ�{ ��թ���{��a��e�H���7�F~�y�(����1o*w��!s���X�#AZP2���5�˩���.|�#`���g�W��g|�Z&�4�mҫ>��?B6��!)�8��AL��+9��ٕ���F8����o���sp%�T�8��~����?�
��`���c|}��BX��w-�!y��Ȑ����,���w
���#V�&�t����'f��z{9k]6L
>N�@tc�ϒ���T)$d�I�v�Oi-*������P�)����w&|���I�����O�2��f�<�R����CX(��_vO�<��f�� ��r}�Wq�F�;5� �a��Nc�<Zl*�g�w�{;*��3O<^e&�e�3������0/SN�f	���!kJ���-nG�S	��P=��`�������1\W,�s�d��{���~܅�ݞ����P,2B���4�����,bWX��s�x��X���7�&.�R�3ԭj���r������@z�������uŖ6$\K��D�<��0����;
�iE��&r��W�h���p׊}MX�]y�+J9���Y��7|�/�Nv2�A2����j?d��8쒪\ζ*)m��&(e�湤{��&������Y���V�����X��T��~b�ģb=4�W�e� ٦i�� <�E��$[7�/�Ma|6��?	+٪��]^5��I,0�n��w׸[�	�!�`�(i3�J��K�8 ^��q� �o�y!�^��R�8�!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc(#`��Gcp��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�/��r����N{a�9O��^���!u�;�Z��uq9����ea�;y� ����t��X������tS���}n/a�τ,Sp�}�f60k��{U��֜��3��TG���PIÙ=�H%T��GF̧̈́��)�ܐ�ʟ�]�AZ��:I�"_��V����p{���,�#������s�0F�2�^���=���8��/��m�����W���9�uP��@)�|{eqG-}p�!�g�[��V�/��+d��;qVeE���jO$xU]c�h�����v�ј�"��Z鎬�������(���/p���x�CyW�f�tR�wX��q�\E��0� wp�R�4��-��%M�rs�i��UQA$��5�%]���a(􆿳����^��Y&X?r>*�3���f�]�!����M[��Ǣk/�z�xEQN�By3��<�]�!����M[��Ǣ&��s���qN�By3��<�]�!����M[��Ǣ���ꀍN�By3��<�]�!����M[��Ǣ@ E����Yl���#�]�!��	Ǹ�y85�;{��T�|>����n���:<��jq㧵�0������0���S�BgV�0�ם�k��L��]�>q�P ڨ�| c�]h�۟�r�@m��+�ވΦ�籢ֺ�9�W|�.Ҩ�5����`K��GFwk��V�V��D�BzL͊�q��!P�E��S��c���>��4�?�g?_��<'P��!jcCA�T�g�v�'s��k� �$��Xo�ii=���JHn��z�S�Ơ�=���\6��.�E�]��c8?-+eN\A��վ�$��Xo��ڭ���s�b9����9�P�rS�b�8Z���'�e�����"�?;(��j67� ��˽��r��B�����O:�	��kIÙ=�HAmY�f��Ea�8S���e�y�/p���xL��fl���=��fLRJ	zh���$��Xo�8�g^��8���ތ�1��\�v��\Y:����QB:�0�϶ߨ�,R���9�"�5[�=�5x�џ�1�?"�E����FZ鎬�������(���l
��������ӯIJ ��`y����@����gG<x�uz���s��um��Q]� _�rs�i�_n����B�Pcsù��L;Л��|#9���b!��u፬!#��Rh�5בvk!7s�9���o��S8�9���SN��'6���;8=�g��U-�e,%�0g���[�=�5x�k�A#�G=���-�>�Z鎬�������(������oD��;mQ��8���/����,D��{r81�lMȆs�򕲠�+�J��Y�{'%s�rOw���é#7ۏs|�Q��Y����2����..W���ۗ���WYHp �:�Z��p�]�!��	Ǹ�y85�����S��C\	��K(����`y����@����gG�������E3-	����V���˺�rs�i�_n����B�Pcsù��Q��Y��ټ*w2�562�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���́�	[��x��;���m���ȱc��/�hz�W)*��!km�����P���L5ӥ����׼��N� ����<n��#Y��"�E��h'�|�W#��P�!͡=5�n�NQa"_�	Z�6㑤3���S� �_a�?=t�ܧ�V=q��Rȡnrj��Gowx.�=i��yU\q��+��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���6��W� X��V�+�3q�bx�#�;� L5ӥ����S�ۗ����f��DE3-	����o�?{/T{9��#.���G}�j�d�t%>^�ߦ��|R%��<��0n|�!h�b���t�m�+�L�w�s+�¤]�o"�s�8��cEp	���>P�2-i_q?�y��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc#��x�y2��5"N�W��\~F}-�=�"��n���Z��G�����M���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�`<Y��spx �M=�#�`<Y��spl
��������ӯIJ ��`y����T֣[\5'b�8�jx�WaU�EKn�+D���ہ��!�#7ۏs|�L;Л�����V�M�$� %7� �@��&}��}j�=��Y�$��J�ֶ�7r��;mQ��8���/�KZ	��\#����̵?ov{��lw	�X�I;���
��vK�Po�Q�>°�������F��#�k�i���A߹.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�����47��.��zN�_�94��"-t"wdC���ѭ��Km4rz��s�8KT�6?���M��,:�-���F����D���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ˮ4T�G��c�{�#�I����~uZ鎬�������(����.��$�ʝ.�&J�!-B=�6f��Z:S����b�Bϱ�O�E�l`8x뛀�������Z}�Y&X?r>幛o1����k$ !�`�(i3!�`�(i3�]�!��	Ǹ�y85��X��I�ՠ�;-�]�`<Y��sp�¨�M.c4AԢ�a\�T��}��w�x�z�2��=�A������h)R�Rl��&k@C�Ɨ0z�cUL��ddՅ<T]v1�_ُ�T�'Y��Y��{&���'6���;8=� ��g�SEս�9�j�[O�x��Q!�`�(i3!�`�(i3!�`�(i3!�`�(i3�uz�#-]iL�1p/-�����̵?o����oD�d5z�R��5 �8��B��;,����ӆ�[W{b ���Ӧ�ȔA
i�eL!�`�(i3!�`�(i3�#�-�p�Y�{'%s��$��S���b�Bϱ�!-B=�6f<Q�vn��l����I�/=k��T�'Y���`chT�!�`�(i3!�`�(i3!�`�(i3!�`�(i3h큈��]v1�_ُ%�W�%�KY��{&���'6���;8=� ��g�SE���̵?oJ�
�����WYHp(�e�	�<���!���c�A�L'�ɻ�L�1p/-��ս�9�j�����oD�d5z�R��5 �8��B�;j!%�)��=���!�`�(i3!�`�(i3!�`�(i3!�`�(i3P"G�wk�Z�d-�~Ee�1���1�����b��[� p�!#��Rh���K�6���!�`�(i3!�`�(i3!�`�(i3!�`�(i3�(]:�z�-ﱳ$�i���		Aqf1�.��N����k$ !�`�(i3!�`�(i3�]�!��	Ǹ�y85��X��I�ՠ���aٔ^?��[+��.Ȉ�;1�˚�!��JlR�`<Y��spW9��8V���ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3AԢ�a\����R�?�������|Pcsù�u�ȭ�>ѯN��S����Ra!�`�(i3!�`�(i3!�`�(i3!�`�(i3-{�+2�p6�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-����&T�ͪ͌�R�hb�,�#N�Trm�l$v��:�_���
�LO��#l7y��6�����}7�
t@Uٻ��
W�,�Y*��h�e���P2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���X`
�2�y��|JS%_���@g�6�o8:4�I���c�90�Ǘa��x���+�^n=\f�5>�|��wLT�z���5|��7�癆cgQw�c4~Nr_�mS8<�n!�`�(i3!�`�(i3}�gv�oE�[��s�A>�xw'��M�v�����FK��|�H��4"{k�h�+]c�)�dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(�8�u?��I���?B��#Ɵe�*|�÷�Wе ;�jmT�#��"����G��Hb� h�ҩ����"sS<ACd�\��l
�����΃0�d]ZM?��y�!�`�(i3D�wP�/�w �%�|0�*b��93�|���1+$!�P{� ܄��w�ƃ
ᾆ�x�T�\ ���:5A��p��w�w:�!�`�(i3D�wP�/�w �%�|0�*b��93�U���c�!�P{� ܄��w�ƃ
ᾆ�x�T�\ ���:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx|��wLT�z���5|��I~m��DL~΄gO�3��|��[�侰j���