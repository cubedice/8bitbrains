��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��]	h8��`��(	�t��L|�w.j��6��H4ي��2_)��:B!�b�ؐ:�{T�{df�r�<�XD�* O�:�k��X�.��ѫ�� �mD�?ea�8���`8��xS��������]��;�I�����)O��Ξ4�"�\�� ���K�O�{����a�s�O�ET?�(�c\֣�I��B���t��|U|�/֚�?d��Y�Y0V�MG��U�;�\����vg������W�aeYgA���z�Ś��
��H,7f�t�뾌��lr�)OI3��(�!����Y�f��a�Z��V���a�\�nq�M�4�Tڢ�]���b��в0FXt�����G����a�����(�I�?g�f��u�H(�3$�����$.:&R�nU���T�����\�4�sW c`k��Zk ��U�i��-a�<�*:>�~�MUs ˙=�=���f���e(�܀Q�ӎ'�d0�(""J7�1��%��.-4����] '�bJ�~C�an��N0r�O��C��0��$�>��w�SA`�/T-B�}8���u���;�'�� +�ۛ���p<�������,�\�H���UDcKE#�4*��1���l�,=�2\��c�鿷ŷ�z����~��M�{�ڌ�2¾'�UB�m}����������uS �����t=�L��^E�h/�����a畹�{�ڌ�2���-���t�VK4��i�;�t�!�k]�r�r����SU8")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[n�+�Uz�QL�W*g;Xv-~x��䂁!�o��c��(r���U�2�C�b��}SO,F=d9�[l�&��q�©���H��JnXe�+�Uz�QL�W*g;X^ �Y�)��H*�m���b��y�.V&��B֥�(����5�:n�|����Z=%�y�g�M)ԉ���S����j�}�I/��=��K�R�/ؒ^�XzL͊�q��UG�s�����v��z�N��������\�v�X�zgq����2��̪U��֜��3�b9���j}8o{:�����Y�V�����ϲ�`�����"IÙ=�H<z,Ҽ&W����vcy���n����\�vŢ+���I��]V�H7'�5�}�]��Ϟ��D	��U�l>o��|�`��-���؍��R��j�.(Wx*��|��pe���b������5	���]���>����C�h�'f R!�`�(i3��|g�Y�'���Xw�E�i�m}6�B�r���E����F��j��\w��0]EOJ�uxm�3���w�@V�"�����/�]�!��M8���	D%��_�ͅ��/��=��K�q�?l�_��ct�:��RE��W��_�ړ8���/��^����r��H�+k&v�Iz��j���'b�t	�U���C��O]r�<Uee�,�Aٺ�H�NI�:7�N�5�%]���a(􆿳����^��+��%�k<�6��w������
L'���Xw s4S�'�i��`�z��GZ>.�0����[���׿j�h�<��CyW�f�t<|����faՊJ�e:[e��mea�8���`8��xS�������Wa�b����y�E�nwE��S��}|��XH�����,>$+W��� j�(����5�:n�|����Z=%�y�g�M)Է\D-�۪�#�h��/`�㎏qló��|����=%+]Bo�A;h�F��O�i���Z鎬�������(���`$�P.eE���lC��U�T�\ ��y�.�`L�H��WOg�Tܔp�l
d�o�R�GI$��ǂcY�~�s<��MR�������c�A�L'G~��6�7�5�%]���a(􆿳��?ƾ����� R�B���B��㎏qló��|����=%+]Bo�A;h�F��O�i���Z鎬�������(�����@��
���lC��U�T�\ ��y�.�`L⯳5����3�ܢ;|�z@��:���GI$��ǂcY�~�s<��MR��G&Tf��@��
���lC��U�T�\ ������q�f@[�=�5x�� �i�#n{Pd�Ӣ8e�2l��4��a��se�ξ������ei4����/��)}���/��r��Hқ[�l\����	N^�U{xN��i>r�<Uee�,�Aٺ�H�L� s�j8[�=�5x��[N�&ѐ��P>Z��e�2����&���Z02��`�z��GZ>.�02�0]�J}�
�?�?KYC'v���NE!/{Pd�Ӣ8e�2l��4��a��se�ξ������ei4����/��)}���/��r��H�"S���X��`�)�	�%{�;����f�kN�ı&l����[}�@��L}�
�?�G.�:��@B!�`�(i3��P>Z��3�ܢ;|�m8^����M��ҹf�f3'bҷ�4K��e�3�x+�@��-��u�Y�KGAc<�p{��K���'��e�V�/,�i7N�_�z*K�/��=��K�9T��,�����Z��y#׬��5�U��)���Y;e�iKI/B޾PԐ#��go`(&�L�xjzӝ���I(͂��-�����2��}�������Ə��.A`��x��nF���<�W�.�P�	��
�Q�}�G�dE�h�����?uA|�d���{_8�Y��=�}�Vݨ��}Dq�f�)�{6�U����$���͜P_�_S:g�RMm�o��'����Tj��^�G�E�BS�+��U�,�P!6���r����܌;���'����u��r���2��}�������Ə��.A`��x ,��rQ�f�6l�}��}Dq�f��G�dE�h�����?uA|�d���u��g��L�}M�9s��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��jr��*�tt��϶C�;��|B *���ۃ��5�Acaw��*ܐb�m��v��z�Naڕ�!�c���Z��q�\E��0�����?Fe��1������Ə�^����r��H�Cw�Hm��mj�B��Vo�I�0hK6j�"Hs��!�2+�*䟭�ab<W��.ʀ8�t�|2;$�JأͽgF"?�Q��ǺΕ�f�f3'_��s�֙Ш��"x���������o��_�Rv�䩲$���dS@Ɵ�od=��¾ȼ;�jmT�#bs��2[�a��o���H�RtV�^��4-�b_X�XV�b�z'hۉ)��d�7�qĹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv���H�����Yu��� ߛ��usȸ�"rR��U��3i�z6��s�u��p��V�M'��w]Pi�#��R!�`�(i3=��,���H̷_��yC��S8�����ZK����t����>3���w�@V-���,W������0�� 7�J�[|�m�ߕ��[���#�!�`�(i3�Y�m�k?j!�`�(i3�/�cLbŪ�����:Y�{'%s��$��S���b�Bϱ��<��>��h�EtC�<�+������L�*dgN;�r��H�?X���V4&v��؄aX�
�:qEp�;�P�t�5!�`�(i37�A��\R��c���鿡�t����>3���w�@V-���,W������0�� 7�J�[|�m�ߕ��:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6���@P?�(w�R���y�sL]~цߒ�a`p�YXm"Ҩ<���v��z�NFX�5�B�ʏ��Z��M^ۋ'��i7N�_�z*K�/��=��K�9T��,�����Z��PlJ�M�=ĥ��!�IX0F�MV�ҁGG�.Mm-;���6}���(&�L�\���F�`yx�>�+X�M?��y�!�`�(i3���_��������صW�my$�N��o�/���;
�:qEptiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3܌;���'����u��r��!�`�(i3�.W��&k@C�Ɨ0z�cUL�����>R�w��뱐�!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2�$�)�vxmiH�f��R�<�t@����,�ǰ����A�z��;_��8W�w��fD���g��3�5��m��� JO��"�5��Dz�͒�p��e"5�O�%E#Pz-j���N�s^�����	}�@�w��˪?�-���ei�^�̷ؠJ��:����{k�h�+&tS�D�'���Xw�j�7����rF��8��E�i�m}66j�"HsXh���(nTVo����6j�"Hs�L*��h��Q���}�x�[������H��<�C�Ar��� ��иܖ��A�.u�r;��|B
y�3~;�>sk8��:���,vQQA�q�m�,�5�%]����8�B���ow_;O
�J��:����EOJ�uxm���#cB;:XSC(�<��>��𱒁�"�ά�o�eHN��R��?�d���&��}V�)c�`�P���w���J���O�������u8q��ǵc��5�%]����8�B���ow_;O
�J��:�����nސ����#cB;,��K�Xmj�B��V𱒁�"�����HN��R��?�d���&�h��R��e�aT��3G?�d���&�[�I�WꐊO�A4ZY�j(&
M�K;��%YM�	�v�3� k�|6�8��:�EB�Z5�O�%E#P�aY��y�`@���!����'d!�y]/�qF5x|���MM
��,=?�d���&�t�{#	�x�jsrCm�k�:��=#��9f2Pih{Ø�F�HN��R��?�d���&�p�T82g�{�Bͳ��;��|B�1�A���^Ta�L �t=-C ��U�