��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��W N��|C��#�N' ���x�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R��
�n�T�+F��W��`h��>��ׯ�=>)m��U���T���딣0&_���X0���2|	p��rw@	@us���)�]&��_	��u|��yq�`݊�|���"rG�
���}�\�bJ(9�{��r�H�����طǪh��p��U>?���>�`\��Yi���u����l�|���j@��"�O��$� ���xI+r�� 0�D�A�f�mXׂ�(ѳsv�`�S��Y�ix�P�Ra����+��a̞w���{ֱ@�W�8d4؇��2O��'HY-�!�5�?�����?9S��m�S� ���������	x]�m�Je{q�Я�mڍ'T����X澗�)�$���:�%�+T%2q򋙔�M-US-�8<�n�У�Ǝ!�ѠV�>!�/�7��u���nEA��x�!ԝ�{��/Ƽ���\�4�s���rH
>TT	q��$�2�����b��ǾI}`�~�MUs �?oQ�%'�s����o���_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3ts�JFAa�ߖ�g��o�4��?����DNZ�j׫���?_W�\I��ఽ��`g�5��!08/?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_E$ô&y���[�nh�/;KYˆz}()pxt4���J4xʆ�7���I���}�����b���q���1�:�Ω�S�T�;Ϗk[�^��_E$ô&y��aC�h�>�N{a�9O��Yk"1/1� =�cw�)&C��4���R$��Ct�z&��ÃlO ܅d^�R@Κ�2���ei����L�IÙ=�HF���m¡;-;*�7��ʐx�?ێ
7�\ZŴ�(??a,����\{F˯�+)�Y-�E�f��Z�>)��p40�zɈT^�`T�W�88�;矷	�gJ�ÃẶ��Ϊ���Jjz�I�~�џ�.���hGD@�F��q���i��I<��fҾ��9��a
�+��8w�=�J�5�o��C!T*Y�{'%s���'����F�r�f�t��6��	���`y������q��ww�=�J�5�o��C!T*Y�{'%s���'����F�r�f�t��6��	���`y����q��G8����<L�|��]���c�A�L'��!�a��5�%]���a(􆿳����^��+��%�k<� -���ݥI��w��,������;�<G��[���ei��"X��[�I�!"lR�^Ƒ����"X��[�d�a�4$�f
�[$��o��C!T*�q���U���d\��N�By3��<Z鎬���������o�	����}��S�)37J*u>����CΊ�?��[�<��z��}�\w��0]�\�LtF��o��C!T*�����2%=dϖ�i�@O�x�7���q�©���$Z�5�8z�E�^�������Wa�b����y�E�nwE��S��}|��XH�����,>$+W��� j�(����5���.�^�9��ǘ^�?�;��XC<�I�$�Q�p�m~|�֛z��8��Ws�Ҍu�����<�սѡ��Cҷ��e4��t-s����eiuKr�'i�dŚ1N��
��D&e�2l��4�y��ɦ�@^7&ģM�&yy��<:�W�_ĵn(���˧�0z�cULjaGkƊ~F˯�+)�"j���b7|#9���b!��u�\.�l����􇃬Tk��A3�(N��㎏qló�Q���l�,�Aٺ�Ha(􆿳��?ƾ��,�&� +J�����|����OxtX+�Yo��Ⓖ���á�~O����}���7�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e���b P_�F����4[٪�E�N;�L���9��Xv7�j��иܖ��A�.u�r]A�S �>{+J�����m���Vή.mH^�+��@}�M�U/��Dkh}Nw��諚��y�[��0���߫�]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�e,%�0g����Ed��>�^);�OA�uW7s�9���o��S8�J�]=��R�^Ƒ����"X��[��Q[R�7����n9읃g9l���z��Q]� _�rs�i�jf� l�Ǜ������CyW�f�tR�wX��}�
�?����om)��%��(��+'���Xw�j�7��ct�:��RE��W��_�ړ8���/����,D�=P��[_kV\�헌k�:A�	S�r��AR1<I�0�f�#/��=��K���ձ�Z��8���/����,D�K��D��`i�m��s�k�:A�	S�r��AR1<I�0�f�#/��=��K��!ҫ0�R�wX��}�
�?�+��%�k<Z it���;;*�}Ւ�~ܔp�l
d
�3�x�. k�|6�8"j���b7���Øf�ƫ�G���N���T	6:��=����זρ5�D��
∺V��܅t�iZ]XF�������́&�Ө��{�V�f��[��iJ�~�Y���(���;����f!�`�(i3�i3<�f�D���X���`>����������o��)�ak�m6"�,�>E��ʆ�In��tT?�7G|`���N�v*$�!�`�(i3�i3<�f�D���X���`����"��5�w�yzw�����+"�,�>E��4];ˍH��!�,���;���2[����|��1�J�a3mPy�S�W�W`!�`�(i3x�]�V���t�����[F�a�+S:H��+܆"BT�(��c����L�{7�ܥ��2�`e7��9��×�>�濖��#�(y"BT�(��c����L�{���D	��U�l>o��|���bǬ�= �zbw��(2�����
�b��{�P}�=]A��O�T=�4e=��-Y�VN�=���Ζ�{QU2����0�5tU���+�J��U<o^.K�}/��<Ӭ�/�"�����_G��?u:�L��Y%T��BP��&��J�UG�s����s�٩���I���Т��^�\7�ܥ��2�`e7��9���I^Ɍ؝�hy�/B/���^!l���Z1����x�'aU<o^.K�}qW8+���?iRPs�&�Ө��{�}+�o�n��iJ�~�Y���(��U��?D��!�`�(i3"�,�>E��ʆ�In��tT?�7G|`~�Y���(�M����H}R!�`�(i3"�,�>E��ʆ�In��tT?�7G|`���N���96!�`�(i3"�,�>E��ʆ�In��t�_�R�Gl�����b���V�Lx{<qH�~�"�,�>E��4];ˍH��\B�����g�q~[{Q�|�\m��Z��N�l�B�r���E����F���8�TPm=_g}b��t�S:H��+܆��K����!�`�(i3зq8�Ј)w�<�_N�-Ł$��Ь>�#�_���}Dq�f��.��Ԕ�]��3a��!�`�(i3���D	��U�l>o��|���bǬ�=l�����2�����
����7
"�,�>E��4];ˍH����TI��Ԫ,щ�"�t� ��O���}���i!�`�(i3���+�J��U<o^.K�}�d	c�b��8���&�r��SQQv�x�����D ML:��Yg6���=�4e=��-"w߻Y��}Dq�f�(����O�^�|n�M�!�`�(i3���D	��U�l>o��|���JLm|��|#HK��@=���b�A������!�`�(i37�ܥ��2�`e7��9��×�>���`�)J*~���f�A�������E����F���8�TP��@E�`�8���&�'�al��pz!�
�W@!�`�(i3=]A��O�T=�4e=��-Y�VN�=���Ζ�{QU2���A������!�`�(i3x�]�V���t�����[F�a�+#�n�%�<�'`ٲ�,�Xʚ@hY%T��BP��&��J�UG�s����s�٩���I����:�Y���зq8�Ј)w�<�_NX�ʟ�3���M&������h�? "a��%}w�dN����+�J��U<o^.K�}qW8+����8���&����uSj��Q�s΁�a�n��=]A��O�T=�4e=��-��~��A��<�6�Q=	�H�Z����Q��nT��Q#>[��b�-W��^[�΍�>!�`�(i3!�`�(i3���+�J��U<o^.K�}5��s� �+U���z�W�F��X�C+�t̷@V�� �!�`�(i3!�`�(i3Y%T��BP��&��J����$�!h�SSB�����m�%��~?H�?���i�jw�jս�������8�TP��k��p�ݹ��}��Z&�lq6�.ʲPdLG���6!�`�(i3!�`�(i37�ܥ��2����*����i��>�`vx��c6�����b(!�`�(i3!�`�(i3"�,�>E��4];ˍH�v��K.Ū�X��oҍvx��c6������|)i��OP���!�`�(i3"�,�>E��4];ˍH�v��K.Ū�X��oҍ�`��rE����ij~�*k`Ë��!�`�(i3"�,�>E��ʆ�In��t�_�R�G��!=.�
kZ)� [��v���Q:�g�a2�-�!�`�(i3x�]�V��w�7qyX����1��H,\ͨ܉p������aUMf�n�Q]�����	!�`�(i37�ܥ��2��fƆ���?|5#�Gm�X:��+��N�C��(4];ˍH�T֟��B�:УWKŃ
.�Ūz�ȣ)[CȪ�U� ���_��z���u�;����2e�5�O֐V���o��k�I#�ā9���8����W�%kԒ�P�K�T�b��M��d��p∺V��܅\4L$ֵ�j�iy[���ҋX����Q��C� ��!�`�(i3!�`�(i3!�`�(i3k��j �%��:wJ~��b{'�t���s�����s|Nb��'1-��B�Noq�ށ �~K[���#<��z��}�z�-~BLI�!�`�(i3!�`�(i3!�`�(i3V����(��N!��qő��{����gFUӮY�E��vNd�)i���
�mN�By3��<Z鎬����a�gN�3c!�`�(i3!�`�(i3!�`�(i3�����U�#�ҒIs{��f��C�'��"�����q��l0q�\E��0j�iy[���ҋX������S8�=	���/lg������T�\ ���KD��}[e��0�U�S{����<�6�Q=$�D5�bY[XҹvXI)�vNd�)i+�0\�NN�By3��<Z鎬�������(���$�~����$^�V]��}1;Z�减l|�*"k���(ӈ��4��S;UA7��I+N����-���q\��Zt%��m&<g+b󆤐=��{l�f|��rs�i���YN�聟�lҟ�,0=]^	�&|#9���� л�.���N���>���n�J�LQ��w�6�5�p����}���S�)37J*uc�A�L'�t�O5u�l�+�	�g��U-�ee�@Rv����my$�N��;� ��b�� л�o���ߞ����>���n
�z��+?i`YS���*';���3�q���Um��#��*y��+�^@��#	Ͼ7�Z#^L�)�4)	���E7��I+��v��q��y�&؏R!׻�p���f
�@"��wҦ�kQW֑��bk<����-�˳k�L��<�6�Q=�w�3����f
�@"��g�����Mgs�4�����DW+'4"��.B�2g>~qA��@����M�P�;�ȓM�Me���섫�So#ȓM�Me��x�2�Hxl�� ޘ_�9��\�'�������>Q��?qr��Kl3��T�Ҹ�MS�B�|��T��tn�+�e��j�3����&Y��V�贅����OD��G͘B./�<ĩ�46�;:���t�b|bQ��� Ǐ˨�g���!G#�<��z��}�<ͧ�:|�"��ӌ�r,�ttT� O���hZ鎬����=���ޒC>ž_�F���^W��kD���4B'�e��n�FM��`��\n$̱~"��>d�c#�'����^W��k�������!�`�(i3!�`�(i3�Ѳ��aS�!-�+_����1�"`��Ę*��7��S��>z��OP�/#�x�+-�+q�!�`�(i3!�`�(i3i`YS�����9Z������?6z�9�ot8��$��.A��+��T��s�٩��um8:8���]�!��5��E0����|e"� 䉇o�M���!O@T'���Xw�����U�VA�ڦ�c4&bݷ�%O�e��n00�8��P6�Y��\���(����A-u��6�0;��ȓM�Me����ΜtȓM�Me��x�2�Hxl�� ޘ_�9��\�'�U�"�����<º#xH�i�é���Vs��nlH�I<�6�Q=�w�3����f
�@"��g�����R��H�O��	�d[��K�pHj�4�\��F���77AƐ^�87��I+�T���B�H��y�&؏R!׻�p���f
�@"tL�^VG����L1�%TԞ}�{J��n��&�P��k<kbm�ѕ����[�|�"u��ӳ��C1��g��U��q�o�u�/ZB�JU��\bE����Kl3��+�I,�S���R����)�&��_���c�.DٖM?�_�9���{l�f|��:2QYeƈ)P<�ܓ�Y竷b��"&�����'�Z鎬����Ĺ#{��ž_�Fȓ'�al��p�M>�I�dB��{l�f|��:2QYeƈ)P<�ܓ�YSƏw0���:ʽ�f0�J.�A�]�!���\B��Vƺ'���g�>k0�ޏ�OEǄ���]�!��	Ǹ�y85��q幊s�?����H�n�f���\�g��U-�ee�@Rv����my$�N��;� ��b�� л���eY�b6=,����hQ���}Q'݀�=��⹌y��o��C!T*Y�{'%sgeߪ�{$�~����$�⹌y�S�UE^����Cҷ��e�ˇ�h����2�[Q	��
�Q�}#�ҒIs{S�>��{A��"�����f��z�� л��Ujc(h�t�%ho����G���r(�:�f,��iQ��e�Z鎬�������(����} "m��^�V]��}Г����ѓ�1���`���A�O
i�c�r׶|�ل�\I��w��,c�A�L'�t�O#��XvU(�8���/�7��I+�:����fSM0.��4;�. ��F����U�e	�K~9Mյ[+8��V5VM�d�}c��%��'MtZ�R�q�\E��0����G誶@~�ܑK!�����+�yƔ��u����L��>���	��z���AZ���d���!i[�t��#��eX�:&���!�`�(i3!�`�(i3���)x�����ő̓Vo���m�#Y���g�!�`�(i3�I����~u�U�pAa��Ms�����x%�n�{��!�`�(i3��������w�MO>�z*K�/��=��K�9T��,�����Z��'S� U�B�\ٿ�6�P6����0�U��)���yk;���6}���iI9�o«IX0F�M�M�Q��#��S����H����Aj��t�35L��$
8��2�ֈe1tSjv��wӨj]h�� yE֩��V��������;q+��%�k<PNm�w�ާ���Cfĉ>99��A0ok��W?�;�끷�Q+��
ņANL�P����<���}Dq�f��q����q!�`�(i3-������ٖ�A$�P�&�2������èV;�jmT�#"��w6�0��ɗ��zi#Y)M���Fe��-����!�`�(i3+�uB;y�� �i��p�>T��O�{ʓ���/ĀI�r���C.�u�X��I�ՠ���7D!��E�<2fsZ��:5A��p�H����Ӥ;�3Pؚ�-����!�`�(i3�2J�4��/ĀI�r���C.�u q��j�J^!�`�(i35��
.ע��x��M!�`�(i3)P6���2��� �;��$3ϟ��7�4��e��� ^C�Đ���%>�rGO�D mWN���%>�rGO�D mWNHN��R���IX0F�M��?���T.�`��ai:�B�:ޗ���::������mIaF��R��#H+�I��)���W�w��fD\Ӽ�gy�A)��/��;��|BK�B�<�t��I%U��_bM+���C����
&h���ٙ���O�Q���*��P�Vr���J��:���鉌tL�<�}}��=�M���w�MO>�z*K�/��=��K�9T��,�����Z��,��G��z�q'&�!�?�P�����;�|��[*���I��:<nl�l�,��G��z!)�M���r��0���u�����%kR��������֢&@��&��$_��f3��"�2VPڢ7���w�E�V{�!�`�(i3���2wG!�S�@�]_LOދ�������y@(8�4�!�`�(i3���-��?s�_{X4t<� ).�xz�\�{<���u*_���X1'1[�?x���"w߻Yf�?ǉ�=K�± ���.]̌�}����q[�Do�9�ݚ�Н�����$G⃕J��2����)ύ^��R�^Ƒ��f�?ǉ�=:��+���y��̨���u�UgF˯�+)��&�C�/��x��&^]?x�v��$wq�����0��E|�,���6%�a¥�����dw�#�ɭAQ�0G�F�r�f�t�Jb�[���e S]#,\ͨ܉p����O,8�ݚ�Н��M?�_�9��@;w�$C,0�?��ʆ�'T���+�n[���/С���?�T!?��vZt%��m&<�,0 ����
�n��E3���?�K?Y��j3�� ��ݽX�Q�L��!�`�(i3��մO��{H��bf�?ǉ�=�s�٩��$�f
%}�YmC,igu��hy��΅���z�Gb��P�!�`�(i3��O�q�̍�Rz(��g�:�B�:�1��?�Āf�?ǉ�=�@�_&�X;p`�G/�'8k��1��?�Āf�?ǉ�=	�6���I)7*{��C��p�-L��y؍��R��I��)���W�w��fD�a�si՝Ӓ>=:9_�aV��	��y��2���,���H%�מM[p|����D5�|�$�* a� k�|6�8yG�$e\X a⣃_B]�m4p`�Xp�T82g��	��#X�1����������Vo[���˚����Z���2��}���/�^��;N�09h\�`��wd�F+��I��)���W�w��fD�?��+�|aT��3G?�d���&�'��G3#u|vӥ{?�VU�簦D�L�x8�̹�y3����&=)X���37�˱�5�ݚ�Н�{�"���ڥ9��[;�h˒�Ӆ��uՇ�OD� �B�S|�P�DM몴PBoTη��~�������
L'���Xw�j�7������}0`a(􆿳��q'�vqng��#:�LH�ҋX�����jƓ�[���Eu ]����b3�'���Xw���\���]~'�H��{l�f|��rs�i��s�٭�`�̳��i;�������T�\ ��׃X�"��⹌y��o��C!T*Y�{'%s�Ǹ2���_�A.��vV�v��g��U-�eVJ:�~�ĬS�V���<��z��}�\w��0]~�ӵ(r7����b3�'���Xw�j�7������}0`a(􆿳��3pCtA 8�����;��]�JڒLy�]q�I���;E�@���=�tK �_"p��W�W��<��W{0`��!�6qK �_"p�{nr���<��W{0`��!�6q��T�Ѓ�Fu�%r�=y�"w߻Yg�����w�-�L��m+)q����h��@:S,���<C���O�G�}�(C#ƀ��=���a��bǬ�=�M^���B!.��@h�^fC��T�z���,}l#�mJ�0�6��������x�&��'�q�BZS[]N���B
��������So-�>�6C�(�HB�O�=��ܒ��Ek��[8{�n�_ �����p��Ss&	�&�
!�`�(i3�ݚ�Н���2�ͥ�lz\�Q��v�r��Rϻt<� ).�x��~\A�أ�g��~�	�7��7�ܥ��2�/��:M/�ա�^�jj��,}	f��J�/`0�����������}�(C#ƀ��=���a��JLm|��(�a��Tk@�0t�bGD@�F��qW��Ґ�Yj:{b6��P'	����t�\7�ܥ��2��yD�0Np�^���17T1���pY�~ȸDz�b9����$�n�����['Ȑ2��;�Q9�	d[�̮�U� ���_j0��.@.k���n��@��P���"5���q�؅��FJ��/��<Ӭ��['Ȑa:�$�77�}�(C#ƀ��=���a��JLm|�V��_�$2���w�"]W��n #�[��0F�s�ݺᣄ�I^Ɍ�|��yf{��������K70y�=`HV7�ܥ��2�/��:M/�CՐ3��F<@�Bcj;�J^��J�Y�"6��O\7�ܥ��2�/��:M/�CՐ3��F<@�Bcj;�J^��J�Y����ߠTq7�ܥ��2�/��:M/�CՐ3��F<�+�����R�:�%��X�B�l�2�vD���?a@!~�X����Ѵ���Z�����q�����P5��٪�N~����=���a��z>�n�S<�6�Q=�b��(��� �5�v��je���Yt	�����\�����!�`�(i3"�,�>E��4];ˍH��\�Mb�mOVy6RTsȸ�"rRY�<�"��@?P�Zv�!�`�(i3!�`�(i3 ���3�ҺIÙ=�H���mL�0ޥ0D���>M�J<0L�J��2���!�`�(i3!�`�(i3l0��F��j �i7�sp>KW℀4٬i�ۑ 55kU��!�`�(i3!�`�(i3!�`�(i3JHn��z��r9�3k��u���f�:X�T�f���y��̨!�`�(i3�E����F���8�TPm=_g}b��7ݲ���!�`�(i3�*���<�Hr�»�>��-U�f��Q��z�n��!�=�4e=��-	i�/B�6��&�elZ�_Hsȸ�"rR�%��ZJTD�l���tL!�`�(i3!�`�(i3 ���3�ҺIÙ=�H�<���͹W�D:���_�A.��W>����!�`�(i3!�`�(i3l0��F��jT�����NM��%�p@�R+��r