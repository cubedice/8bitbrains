��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω������?9X�1�Z�U���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍C95^T��6\Xa��7��Į�N��=i�@x_\q[�@�0�I���j{�N<��;��� B]�pE���	x]̃Dj#^Da����M�$����o��I�绯�t�z����)�,�˛D��w���旴4w�1����h���������$[G��m$�;�`��v��p�㈍x���t�켻�S���c,31�-elwB(�93;2���Zߧl4���0�?�1~�x�c�>j����d��S�W�>��Q�d����t�mR��:�����-��3���7�Jk�b#Ӡe��?�F��&��;�Éi���W:�*c��,v˶�9�ĒTC��0��`�R&.1� 0��]�������yW�u���;���A��j`��'�����`U+n%K)��k��Ǣ���N�y�Yc���;��sD���L��+�Uz�QLQM��S�O?�4�ʗ
� �AH�T�t��3��e��ME
^����c�:���0�F@�4%�u�L�r��3�jT!�K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s��e�IC�_�\�����@J
A��w|�<��y�~/r�I��
����&�ɬ� VU+I���ť1k�`�tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"���`���l��KJ(𬍝��;{g�P�r�|Aڙ���M�	g�yߓ����<�m��+��$|��;D���J7"���`���ld��q�G�+��T����oGo�Z�������--�p�,Xy�g�M)ԉ���S��(�B4�rs�F�r�f�t?�1J&�|D�e�!��L�D��6S�]V�H7'�R�^Ƒ�ӥ�e%)>�Z��&��J��Vǃ���O�4ۤ�`�	��B�f�\�kA�/����<.+6J!�t���\�Ws��l=�L؅��FJ��G��k���؍��R��j�.(Wx*9��?xs���}�ڍ������5	��]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�e�,���6+�^�9.�JQ!�`�(i3��{l�f|��rs�i�� ��*b��0��E|�,�CyW�f�tR�wX�Ռꢤ�Og�?�e����]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+��A�y�0� 7G#+�Ǘ0z�cULjaGkƊ~F˯�+)�"j���b7���Øf�XA���BU7Ê7�E�4'���Xw�_�!	�\�����5	��]�!����M[��Ǣۧ2���{�ҋX����>��l%i�-̇i�d�?���{l�f|�ό���.ӳ�
�	?�<7Ê7�E�4'���XwI<��f�@O�x�7���q�©�����<������ӡ�L��]�>-iu�`���`�+N��?���&���#�{�0;�}����\Ҥ�Yk"1/s�\"���a���ܻ�9���$1m
_g��c���C�x��T��=}�ŕ�F&|S���T�\ ��3��h=T���GZ>.�0�mm|�5i���RY��ss2����m�5��C�F�W+`�x�oE&�0�3uH�@�ԗӯ��~���Ƒ���s�Y�{'%s��.|Z���I7��-5��6��	���`y����@����gGK�(SQF^P��:w���@c
�}�
�?�K�\7}�W,�a��zr,/'���Xw�j�7��;-;*�7���W��_�ړ8���/����,DB�m�?�]�0���߫�]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�e,%�0g���[�=�5x��|��C%�7s�9���o��S8�/ #O�)R�^Ƒ����"X��[��Q[R�7����n9�^����I��Q]� _�rs�i�jf� l�Ǜ������CyW�f�tR�wX�՟��@�'�ǮD���i#���� �t]�8�[|���U��k��ϳN'R�7h�����t���G�ɬ�G
��\���.�^,7p�J��PW�����!�`�(i3�����5	��{�OF8F���m¡h�q��d[dͤ���!�`�(i3jݭ�F���p� o��]�=�<���� z!�`�(i3�����5	��{�OF8��'�PD���Wʁ��c)q	��u!�`�(i3x�]�V����:L���2*Q=F��:УWKŃ�6�5�p����Rܖ��c����L�{7�ܥ��2�`e7��9��×�>�棩�!s�;�����)�ak�m6���D	��U�l>o��|���bǬ�='�u�uX]�����)�ak�m6=]A��O�T=�4e=��-Y�VN�=��`
 ֢����e���W��9�JzM���+�J��U<o^.K�}/��<Ӭ�Q'݀�=��&�v�xb��{�P}�зq8�Ј)w�<�_N`E�cvR+��}Dq�f�]|If">��]~'�H�E����F�Z�>)�ώ�~+�ݗ,�ttT�r�pΚ�w]@� W|`f���D	��U�l>o��|��`��	4��=����t��cg3/F�~f������F�)w�<�_NX�ʟ�0
<7���j�G�ɬ�Gl�_`��<-��.�^,7p�J��PW}ݡÝ���!�`�(i3!�`�(i3jݭ�F���p� o��]�7p�J��PW�o#�_T��!�`�(i3!�`�(i3jݭ�F���p� o��]�=�<���XΚ��!�`�(i3!�`�(i3jݭ�F�������a</Sn����e���W�^�|n�M�!�`�(i3x�]�V���M�K�=g�H{g�q�SƏw0���D ML:�,�Xʚ@h"�,�>E��4];ˍH��\B�����g�q~[{Q����!s�;�Rn\�_�B�r���E����F���8�TP��IL;��$��8_�8���&�5�w�yzwz!�
�W@!�`�(i3=]A��O�T=�4e=��-Y�VN�=��</Sn����e���W��]��3a��!�`�(i3x�]�V���t�����[F�a�+�ީ�%��w�*�fBg�!�`�(i3зq8�Ј)w�<�_N��M��+?���C&���J����i��:��2O!j���Xg�d���U<o^.K�}�d	c�b��8���&��Ŷ;�����}���i!�`�(i3=]A��O�T=�4e=��-"w߻Y��}Dq�f��d �S|����7
!�`�(i3���D	��U�l>o��|���bǬ�= �zbw��(2�����
����7
"�,�>E��4];ˍH����TI��Ԫ,щ�"J�a3mPy}���C�!�`�(i3���+�J��U<o^.K�}/��<Ӭ�Q'݀�=��&�v�x���7
!�`�(i37�ܥ��2�`e7��9��×�>�����>[Hs�?����H:e���f���E����F�Z�>)�ώ�~+�ݗ,�ttT�r�pΚ�w]��Ɋ]��E����F���8�TPO������=��Z��( �s�٩���I��������|�зq8�Ј)w�<�_NX�ʟ�3���M&�"b8�Zv�l���]cK�Q0����+�J��U<o^.K�}���]�p?ȓM�Me���ta�?Ji�@���g��������"D�
�	+/O�Q� !�`�(i3!�`�(i3зq8�Ј)w�<�_Ns)���'�j����Ja|�~(2"{��o N�{u!��}!�`�(i3!�`�(i3�E����F�Z�>)���0��w�wbk�$+��m�yo���|��Mb��y9xOI���S4];ˍH�'N2��D����&�Q(�6k�4d�k�G�E��`�4,�pI�!�`�(i3!�`�(i3���D	��U�l>o��|�w��Y�ڪE�9�ؕ	�-��K!�`�(i3!�`�(i3!�`�(i3x�]�V����:L����(���E�9�ؕ.R���(>?C�e4-&!�`�(i3!�`�(i3x�]�V����:L����(����&d,4���ʽ��Q\w��B���!�`�(i3!�`�(i3jݭ�F�������a�t����}�(�
4��c��^�
E��#	����J!�`�(i37�ܥ��2��
[���p6I�%�.�p����nZ\�j��fxj�9�t�.܉giIE�!�`�(i3���D	��U�l>o��|�e��A�?S7�8�8�``�ǆ�x�]�V��v��K.Ū�X��oҍ(��.��}T���؅��FJ��S0�:�l���\Kd�!%=dϖ�i�&���[� 7��U-����`kv# �	{��� л��;Tl5�����E��~@�k��ϳN'q�ށ �~do���;
U<��z��}�z�-~BLI�!�`�(i3!�`�(i3!�`�(i3V����(��N!�$�D5�bY[0!o�`ƛ��*Z�h�TD��L��`
 ֢���Ӎ�g�cޢ�{l�f|�t�K��0�!�`�(i3!�`�(i3!�`�(i3�;C@����3a�LD�P�섫�So#�rDB\��1P��#K�SM0.��_��܂������5	��]�!����58*�!�`�(i3!�`�(i3!�`�(i3���@�k�r�;`�L(2��>|Nb��'1-��B�No?V��j�c���yQ2J<��z��}�0z�cUL��լ[po��'N�*	�g��U-�eq����9�K7͍��ճ��)�ȓM�Me����Μt�[�}��|SM0.��ʸ=�Z������5	��]�!��	Ǹ�y85���`*uӋ�n�_����Cҷ��eq(����b�z'hۉ)[텡#����Mei|���-�S��Oy����������n[���/�o��C!T*Y�{'%s��F����0@�pgd@^�V]��}R�wX��<�6�Q=$�D5�bY[�����-VL�q��l0|�\m����(���ҋX������S8�=	���/�cv���٬a(􆿳�tP"7��%e��0�U�S{����<�6�Q=�qő��{�����-VL�f��z�� л����O֮�
�W!u���-����UY֭���F�eO�V2y/��S:�cN���dt�{�Y�Mei|��Ja#���a�7�%��S�ғ���X��4tΘl\	�����:�!�uM������i��T�ȓM�Me���T��G���X��4tΘIy�����OyQ���ؐ�d�r���H��O�	�v�,,�kQ���t�b|bQ��� Ǐ˨�g��F�d������U�We��ǳ̨����2c�8�4��&Y��V��CE����r�գ���VRj8�@ʚ��X�a;���T�ҿ"`�7e�ӳ��C1��g��U��q�o�u�/ZB�JU��Q��?qr��Kl3��T�Ҹ��x���-�z%8;����v{:��h���#6q㢝{l�f|��:2QYeƈ״$(�>g�Y��j3����lj�]�!��5��E0�ƺ'���g�OP�/#�xΨ�	�ǳ��'�Z��똣w�ٽv�yq�`0�|(O��"��"�T�>�OP�/#�x;��C9I�!�`�(i3!�`�(i3i`YS�����9Z������?6z�9�ot8��$��.A��+��U�U~�}];�SS�΅���!�`�(i3!�`�(i3�� л��У��a�p�탯;\߰ �Ye�]r��8���ҿ"`�7e�,�ttT�<6(�S�)37J*u�,�JL����?D�8����9K��r|��8	(1!Z鎬����=���ޒC>ž_�F���gz=��qװ�U�3�?J�J�D�k�7 �:�BF�!���q�%��Ro�����:,:��F�d����"'l��*גǳ̨����2c�8�4��&Y��V��h��)��X'}���.���� z;x���d��P�;�ȓM�Me���T��G���X��4tΘIy����ߗ��L1�%TԞ}�{J��n��&�P��k<kbm�ѕ����[�|�"u���Mei|�J�8#O)a�7�%��S�ғ���X��4tΘ���VC0�����i�é�I���z�S�*��iMOPԙza��5N�ʡV�l��� л�G/1avQ�e�b�����,��Z?m��`�������VRj8�@��"�VGN�Ar��$x(p�Kvv�77AƐ^�8�o�@h�H�o��C!T*p�VU��Jm�QA�Q* r�VU���?��K�U��]�!���\B��Vƺ'���g�J�a3mPy��9����o��C!T*p�VU��Jm�QA�Q* Zt%��m&<;p������l�r��S�)37J*u�,�JL���毘3)�:֚S��~��N���^�S�)37J*uc�A�L'�i����
��8���1�pp���aa(􆿳�tP"7��%e��0�U�S{����<�6�Q=$�D5�bY[�q��7-]P2<WV��
i�c�r�(����O�����b3�'���Xw�j�7���R�|E���(����O��J�[r��-�8���/�l|�*"k���(ӈ��4��S;UA7��I+��$����^�����m�z��+��ݘ<�6�Q= 4'���G0>w��Bw�B�"p�l~z��l$c�� ��e���]�!��	Ǹ�y85���`*u�����7����`y���#�ҒIs{:�Q7?�G�vNd�)i}#vZ����@IE�U����S8�=	���/|2��#�	�T�\ ��^���[B�I��"�^�GeY�]1�
f5��h�1w�0\�o�8�@I��èV!�����+����l�`1M<���8���L��>���	��z���AZ���d���!i[�t��#��eX�:&���!�`�(i3!�`�(i3!�`�(i3!�`�(i3���)x�����ő̓Vo���m�#Y���g�!�`�(i3!�`�(i3!�`�(i3�I����~u�U�pAa�Ќꢤ�Og�[�Qه�o!�`�(i3!�`�(i3!�`�(i3!�`�(i3�MC@����l�����M�Q��#�?f�̗���\�rҖ�A$�P�?�#	*]]�iI9�o«IX0F�M�M�Q��#��S�����,8?<�%�z�-uͺ�s�η3G��Hb� h�ҩ�{k�h�+!�`�(i3!�`�(i3!�`�(i3!�`�(i3A����2�2�g9l���z��}Dq�f��5ߧE4��HN��R���IX0F�M�M�Q��#�?f�̗bV�Y��� v��ɿ���!�`�(i3���t�T�V�r��}�������y�(����<mϝ�j
������h��`�����y_�mS8<�n�ݚ�Н��V.��(�t����BQ�!�`�(i3!�`�(i3!�`�(i3W���y�N�sf�e�}s�dKa���z%t��#-);�OA�uW�H���~���H����Ӥ;�3Pؚ�-����!�`�(i3�L�s;SF`R�"�ѧ!�`�(i36�&��=�K�o���,);�OA�uW^����^����I��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M��?���T��;_��8W�w��fD!�����+t�.�Ҝ� ��(ʧ�q8h�G[�� P��#��s�'	�?��[��羹�.������S��?�F�^C��}��,\ަ�It��+g[����Js�dU�p�[��HFzf+b[w�Qt
����+g#>��?�Ho2����q��3[�T��s���rRV��E���ci�n~�c?D��Bn�W����&!���"w߻Yf�?ǉ�=��4tBu6�]���~��\��,&߰��U��f�?ǉ�=����$G⃕J��2����u~xgA���������6%�a��x��&^����V�͖�X;p`�ct�:��RE3z%�u�܆N����p$Z�"�՗&8�,�I���Ut�es��O!�`�(i3�nxL�J}�U���^��9R�^Ƒ���ݚ�Н�LZ�2e�?k��,�:�N�*�x竷b��"&�ڶ|e���@;w�$C,0�?���Zt%��m&<g+b󆤐=�X;p`�Z鎬�������(������P`��B7Ԅ���6�5�p������fLZ4��s�H��rs�i�H�~ȵ�7�*T�(d�ˀ!�`�(i3�-���k\�&8�,��Q�L���B�'��a��IRZ���Q�L���B�'��a�6+W��-��{����"��hy�^>�����g�Hn7�(��wӨj]h�u��߹c��-��\cZ��2�!�`�(i3�%]�N���&8�,���AF-�ݚ�Н�U�A����!�`�(i3�V��9/���ǖ�!��;_��8W�w��fD� ��(ʒ��(�'�@��x��gwD����c�̗X6ڭ��W�XL�k��]�����aR�����5?�SLq�N��	�<���|1I&��ڥ9��[���"��Y��uՇ�O����ݭ17G#+�Ǘ0z�cUL��Jv(K�V��1�.ΈГ8���/����QjG������'�Z鎬����r�V8>���o4Î87V<��z��}�\w��0]jC�p�����N���^�S�)37J*uc�A�L'����f�.`�G�	����6.R�wX�լ��h�3dn�n��r�ҋX������S8��y�)xʔ�ɘ �V�	ᑭ1�K����`y����1b�"�����!��� ��]�!���Y���f,�r@h�?I<��z��}�0z�cUL��Jv(K�V��1�.ΈГ8���/��� ���D�]Z�Vy����S��#��̻�Yi#���S�U���9Ҥ+��o��s4k�r�j�b#�S�U���9Ҥ+������p���r�j�b#�S�U���k�_�|�ɹ��I�"&`�A
�M^���B1��?t7u�`'s^�`}��AyEy�5`P�~�?s�_{X4x�]�V�����TI���0D�Ub��5�%u�%r�=y�"w߻Yf�?ǉ�=�F9�^ӽ?�Y0�
n7A��^⠻rRV�����K"#oս?�Y0�
��аJ@o�C���j#��|_w���d��G�P?s�_{X4t<� ).�xy<�@=%�m�ڨ�hծ���aR�Q�>σwE����4������y�;���g��d�6��mo�C$�:�;��K:SGD@�F��q`E�cvR+J]���q���>�SS�]�/v�]�9m��� ��
x�]�V���\B������������_v����4�F����>���=���a��z>�n�S�(�a��T��պ�}�GD@�F��q`�U����uEe�t�/Yi��}Gz�SVL��˚�'n�^0o���Zф��t��o�51��?t77�ܥ��2���C�0��(���������l������|�7����s�ݺᣄ#��̳Իt��o�5!.��@h�^x�]�V���\B�������������`
^8�J#w���`�._��4];ˍH�O������=���I�Z|���勤U�@k����c�)0#GD@�F��qX�ʟ�H�Ѱ,���e���}��+�'��r��Zw|�pMGD@�F��qX�ʟ�H�Ѱ,���e���}��+�'��r��)0#GD@�F��qX�ʟ�H�Ѱ,���pV�����ٙ�����\�}��n�4];ˍH�T֟��Bg���j9�0��_o8�
��Člx�]�V��v��K.ŪQ�XT�~R��/�dsE�#o�C"Jżsȸ�"rR�����P5�D������o!�� U��!�`�(i3���+�J��U<o^.K�}��2���֩��)�IA��y����U�����bWz�>H
#Ћ�!�`�(i3!�`�(i3�b9���:&�>��s�� �5�v�^*?�z�̒�W��:�T�!�`�(i3!�`�(i3"�,�>E����\�v��_�R�G���Fz�Y�b>bb�v��UP�!�`�(i3!�`�(i3�Q�^�y�zL͊�q���?�-���!�`�(i3�i(���� w���s!�`�(i3!�`�(i3=]A��O�T=�4e=��-"w߻YKW℀4ٵ���d�|���=�Ҹ�S��F��u2�k������U<W�L�x�]�V���n:�t�c{DJX</���m}�ɺ5w��X�N����p$`�̳��i;*7|Jr|�!�`�(i3!�`�(i3�b9����4�6�tڣ� �5�vž�x��&^ɘ �V�	������#!�`�(i3"�,�>E����\�v�[�w�������aR�?W��;�