��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��:%��Z���xN��g�.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I+ĂiW,���D�+y[ف���rn��mo����/~.)��3�(����C�X��2�k(����)O��Ξ4�"�\�� ���K�O�{����a�s�O�ET?�(�c\֣�I��B���t��|U|�/֚�?d��Y�Y0V�MG��U�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|/~.)��3�(����C�X��2�k(Qg�@zh�S҆�|n������}�K�~^T�ɴ��b��9J�Й�m�z\H�� 0��~����p�:�C��JS�Ȕ*Ĥf���J�D{g�P�r�|AڊR$�޵�y�͌�4r�O��C��0��`�R&.1�s߬����M�!�֓��u���;����\_�MX�9�I�[��On�AN�.5f$��F�Ŋ�����}�K{ɈC`N�z����le�kI��Ř�^~tҦ,��_!���5�NnZsA���r�O��C��0���/���k���_0��*�Ε�u���;��.~�Gj'��w9����`e�TS�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l����2�C�b��}W�����%3?���kW���;��sD���L��+�Uz�QL<(�P[H��Z˻r����I�?g�f�L#����2=�l����2�C�b��}�@���,������0�ea�8����:%��Z��vDY�όW�_42K�,\ަ�It�k\,آ()���;��G���9��'n�^0o_
-��[�����Kp&�@���k��l0��F��jT�����Nb�?49�����_�\G��4�	B45k�c��`��'n�^0o�!���!��x�	�2��g�P�e�9�:�]�^��'n�^0oM�D�;��-+0�l�R<�q��f�}��Gظ0���������5	���]���>����C�h�'f R�����5	���]���>����Cοƿ�d��������5	���]���>����C�?KYC'v�������|g�Y�'���Xw s4S�'�i��`�z&"hkIH*���>RTت�I7��-5��6��	���`y����ꢤ�Og�[N�&ѐ��(�
t��Y�{'%s���'���ը��_�\G��4�	B45��lC��U�T�\ ��Tǯ�!�tӱ1R�m��+ r���7���?�_�N��;
�'�����N<���d�k��Yu>�G Oag�qod�֓��+��T�����h�6ؖ�(����C-C:����-;���:vޫ��%�%����=�ܔp�l
d�o�R�GI$��ǂcY�~�s<��MR�������c�A�L'��!�a��5�%]���a(􆿳���2����.��DP֞ �����Ə�i�w!Ŷ���=�ܔp�l
d�R�.��On��M��Ґ�m��[��^�7��u"�$��Xo�����}��!�z��$�'��C0�$i��k��L[���Q�Lmb'}-����C??`J�X��9cѶ�^���4"��"}�`�W��f�(d0iV�6IWJE�\��[�B�9Cd���*�=��X�<�Fk R- ��-��; &+W���F�^�Y�7#�xI��W��_�ړ8���/����RY���+����JT؛>�a�W+`�x�oF�/iu��+W���F�^�g�&�0m�H?�Q�q��ʃ���_����,D�푧)��΁�a�n��v��*ࢢ�2ا@���Ч�O��R��m�]�� �k'{B����ݳ�B��~� gWVbT+踫g(�r��3c���jj�#W�U��ظ�d���!i!q��V���A��u������<"�`�it]v1�_ُ�����Ə�r�����]+W���F�^�Y�7#�xI�~��;�,w�R���y���,!���BȀ����&M����*�Jͱ�F�a�R8[V��M*C.H���{ �=�%�H9?�l0���d���!i� ��鶯bu���Lo�u�Y�KGl+r���%iۋr(���w�Ε<ÚP��h��d���!iO.C�+��uK[F"O���%��ɶCmsW�C��y֘������Tؿ ��Q��d)�I|"nC"��:�%iۋr(���w�ΕG��Shh&5�O�%E#PZt%��m&<�e}�æ���o��_�Rv�䩲$���dS@Ɵ�o��6}���iI9�o��ݚ�Н����"sS<�0�zG�������&G!�`�(i3!q��V�ys��e�sb_X�XV�b�z'hۉ)��d�7�q�!�`�(i3�Ro�G/]%�z�-uͺ�s�η3G��Hb+�����;y��v��\���
^�ݚ�Н��H�����Yu�������&G!�`�(i3SƏw0��A��6��
�g�����;�7��w�@z�צ�,>�����BHS�/����OY'���}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3��ܐ�}�|�:���	��C�Y�\�w�R���y�U��\JD�GLPP?����.J7h����8�ϋ󈷛�'�%њv�>钙���{�v�(��@��$r�f>x�:	�W+��W���f��p��r�d��{��A$�P������5d�`UNP�C>��Ӛ<lȕx�!�`�(i3�r$ɓǃl[�Ƶ�1tSjv�!�`�(i3��hY-N�g	'�^�#u��nF���<�W�.�P�	��
�Q�}՝� s�#04~B3��������h��`�����y_�mS8<�n���F�P�7��S��h��d\�!�`�(i3�
�t��T&���LQ�/81tSjv�!�`�(i3!q��V�ys��e�s֑�3��/������Y�x���|8�ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5
�:qEp$�)�vx�ܛ�Z���}Dq�f�����,�ǰ?%{B��0B�t�A���I��)���W�w��fDe��f�ۚ���;_��8W�w��fD�9V	���8�DKIͰ���@Z���rs�i��r������(&&������it	�T���-M+��00�tO,���6�6����D5�|أͽgF"?�Q��ǺΕ��m��[���^�̷ؠJ��:����}V�)c�`j�Txk^�ԡ�/$a��F˯�+)�+#c����nS�3�ǻ��d���!i?V��j�c���W�gD������?KYC'v�����$�/�x��HN��R��?�d���&��}V�)c�`aT��3G?�d���&�[�I�W��w����|�7����c