��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVD�6�����;��sD���L��+�Uz�QL�]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUP���*+�[��������-�7�5��;��sD���L��+�Uz�QL�]��;�I�����)O��Ξ4�"�\�� ���K�O�{����a�s�O�ET?�(�c\֣�I��B���t��|U|�/֚�?d��Y�Y0V�MG��U�;�\����vg������W�aeYgA���z�Ś��
��H,7f�t�뾌��lr�)OI3��(�!����Y�f��a�Z��Vv�c
���������
&�[��%Fc�;B�@����wx0�<�·�
f��o ��v����qB/�&��w~��19σ\���F����92@�+���aA�O�_��xz8���"�^
 B]�pE�er���{g�P�r�|Aڙ���M7\F���r��RL�a)�Vu~c!��,�%���)0!�Xl�!��5]�H�u���;�;N��;�DnAI���^t�5'KL[��I��'��jT!�u��w)�S�3k:�(�-7��Mv�9*���f��^��#ߪ8�:r&@��=��?��ذ��8")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcl7�Fmi�E+���WY`�`��yXi9�
�ѹaB��Q�/,f$�7Q0- ��Ck�fÜ�2/�r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[n�+�Uz�QL�W*g;X~09h�i��I�?g�f�$��P�xZq��t�1�:�Ω��
�/�r}|��ι%9��oGo�Z�J��ݪ���AOge��L7���%U�"sj� �<{g�P�r�|AڊR$��^[����CԞo�$C�I7��-5+Yi=��o�IÙ=�Hr<�Gf��p�m~|�ֳ(��	�4���ތ�1��\�vņ�Q�]��7��k'�w���j����r k�|6�8Ln��S�W�mV��5f* &�a+�p�m~|�֚?��]t��G�p�P�^[_�e��IÙ=�H@���N�)�I��'��3
�v�v-}�	mpǐ�=�一IÙ=�H��
#�_�I��'�nQ�rV�?.��	޼�\�v���GAџV�$��Xo��Q��F����p�X��#�ڊ<?@��[	J��;hΕ���ivc�f���2�خa�>����n8���ٳ��溂�U~܎VV��5����`KEfVNNKi0j@$��U� ���_�ĕ|G���7��k'�w�W���@y1*T����)w�<�_N �VL�(\-�J~׶�7��k'�w���j����rx�y�Zgl����ܼ���\�v�T?�7G|`�$��Xo���~��1�51	�<�����ȳ�%�MZẶ��Ϊ���Jjz�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}��z�C�f�9��/jC��Mw���1�Z���=�Ln��S�W#w���	(���B���Q��ǺΕR��ӟ-�!|�α+�5����`K��x�壃EE��W��±�sR�{F;�f��X��Ye�?����5����`KI�J��#Kl�Y�7#�xI���|�r�HzL͊�q��n�/��}�������g�{�]4�W/S��8(�E���Kt�+Yi=��o�IÙ=�H)��\a��R���w(��ES���v�8:z�ED}���w�K�̄�Bq��f�� ��~m*�S%���^̽1��H����8�A)�V��/7��k'�w����T�ɑk��!a�tc�&ck��1#��Z�����XP��Ȍ�`�>�fr��VYW\-@��F~*7���&�_���/���l[{{N���zL͊�q��]��B���
_g��c���j����rN�ǁ�f�TJؓ���!��\�v�n��l���z�@ʶ��o��ۜt�[e%ސc�g;�C�2�8�aq��@�)d�8��;���N�i���
ON���:�hΕ���iv��b�7�*�7`����M�Z���	�b9������E\������Q�bI��'��b��v݋N��������q5��wb�S��V��\������� ����;*��k��J���\��иܖ���(��K�K)x�?{���x.�Knq�I��(��f�� �:��#"�RҔV�w�Eh�$��Xo�;��7�"� ӫ/��mk�79�����\�v�ʋ Z4.���A���ۖ)t���sCJ�	�LÆ�Ǒh�~���;
l�ć5����`K��fx'v�ao.\C�k�ף�D�~|�^��
�>IÙ=�H!f+`?>gh�5����`K��M���o�G�m�??2{���zL͊�q��n������I4��欱���j�����ճ�|9O<9�Sz����M����A�m�(���.�Ub!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л���U��u��Y��)�>����
|�NwWk�|��{�ru�?�=�r�@^7&ģM�'n�^0o�<:�W�_�l�J;�Rg��dT�W/S��8(�E���Kt����ӯIJ ��`y���]���.�#�.ZVRѿUJC���d��)Dq^)_R@^7&ģM�'n�^0o�<:�W�_�l�J;�Rg��dT�W/S��8(�E���Kt㲎�������°������R�wX��
|�NwWk��
��D&��:mӖ�|�����V��ߝD9�{��灊�O�i��Ԓ:/��N��I7��-5���ӯIJ ��`y���]���.�#�k�:A�	S�r��AR1<�N�؆�B��W+`�x�o���{��&�e�5
��Ib����rs�i�jf� l�Ǜ�����°������R�wX�ՎF���הtzy�g���+����q���M�I�h��C��-��JHn��z�Lqܳ<��J*�Rs�0䁛����$+�w]�B׿�ġ��,����m��E��T�
���A.o�G�m�?[���S��IÙ=�H��"~6���aq��N�SY����#���F"��5��h+�$��Xo��I;��?�;-;*�7�����|�r�HzL͊�q��C.W26K�~�J�� m�������.��R�}vJ^A"�=�f!��$��Xo��I;��?�C��[�����I���'����=���aw��Y�ڪ���Eck[�x�X��u�?�=�r�@^7&ģM�'n�^0o�<:�W�_�l�J;�RQ�y�� Y{q����'6���;8=�g��U-�eI\�53�f؀qjZ��H@H�֦g�㎏qló��|�����V��ߝD9�{��灊�O�i���Z鎬�������(���o���ia�ƃ
ᾆ�x�T�\ ���( ���S�]��i�"�;���[���ht[�����N:��,��g�7�s<��MR?,��l����>�	M��}�|�݌�˅������� ���9��c^Ǘ/�;Ʉ��W|�M��	�(̲���-�t,�?j����y�N������b=��l�p��i��L��\���c�i�w�Ah*g2��m �A?��V �-��7$2ӔJ�V�	l�JHn��z��p�Sg�3 ���t��h�/a����C4�O+�j~hx���C%�"�uI��'�ct�:��RE�QS����>�b9���S�nU�&u������I��(�G�̅bGc r�p͟�kn@}����5����`K��M���I�m�J�Ln��S�W�
����uK�r�&U������G|M���cݟ�*hjY탌t0�^-��Ys��3�����$7���@e!�}ICq֌B�[v�\��O6�[c����k!�M�Z���	]���.�#�D�of�7���A3�(N��㎏qló��|����=%+]Bo�A;h�F��O�i���Z鎬�������(���`$�P.eE���	fd�L;Л��<��)�A�'�V&����<�#��f2��-�>��)Ȁ!�~��_��r���~3%jA�L�Z�;tm(���)j��q�hY��x�h�@�{d��L�'��d�7[Z�^>L���K�^��x����N�47��Îq4gك8�1��A3�(N��㎏qló�EDF�:�r��VYW\y]/�qF+Yi=��o�IÙ=�Hw¹��<d���	fd��Q�b��3�+���LQ���ƪ���������r�}ٺ�c�ˁD|���xV:�	����4#m�hU��-7��k'�w���j����r�C�M$�1#��Z�����XP���h�5,Wl�/�O'�=�c�r#�_�^@�����8#����%�$�yK��L֨Kc�?�$��Xo�e_�d
���ݪ��1#��Z�����XP��ȗd�uY��K��T��p��`�Q;?�͆�%l9�e\EV	7�j��B�5����`K��M���R'),��`�?2{���zL͊�q��*
�DWo$�}��M�+�C
2��ܗx����c�hm�i�]�׼�a�r��AR1<�N�؆�B��W+`�x�oP��@t�&�e�5
��Ib����rs�i�eB��P�ߘ�)�Iƃ
ᾆ�x�T�\ ��D9������$��Xo����Ǳg�P�e�9��<���h��'n�^0o�'vX[���?� Zh�R6/��������рӚx��	��x���:%��Z���d���F}���3Yc�#�<�R����h�$$����eR�ʨ��_�\G��4�	B450M�/�s���'n�^0oQ������ݪ��A�wd^�۱g�P�e�9��=[��7��k'�w�5kj�Hn�wk���Ln��S�W�bOM�P�C���_�\G��4�	B45�EOs\�̞��>��3
�v�v-}�	mp^�{�c4p�m~|�֙X�D��U9����u�I���'����=���aWc;L�\VW�ȏ�k��a�s+�ҟ�r/�^��D途�؎���ɿJ�:9�2����rR#K�p�k��M����S�	7�i�߸B�9}.�Б��+�B\zm�x�R���-�a3�i�a�>���t��.�Չ_:s�83��˶�D�;K�I��'�U����z~+Yi=��o�IÙ=�HIR*�fN���D>x�N2��m �A?��J�8�+|�.�� �
aK�)�[�Ặ��Ϊ�Q� ~��
|�NwWk�l����4v�7�ZS��|����=%+]Bo�A;h�F��O�i���Z鎬�����׃�Q�.�I��'�!͙��04nԴ�V����U� ���_tE��gVB�3?�J	QT���cP}()pxt4���J4xʆ�7���I���^��p�m~|��w��&�{c��n���|��6)�ш�Ψ��F$��O�&��:�������#W~(�2��yT�n�g�Ӯ�Ⱥ�y�Nb�3�G4R^h$�@Ak���7��k'�w����%iz	�d$^����$^괜�4]�k�1 �O�ok(�o?�De��ӆ� ��U5�\�E�o5��O�/��� �	�q�^!��.�I���'2۶��R���҄��3Z`
���eH5��Òo�j>��i6�0w�mL(��ߠ�����G;M��
����o�4H�/
��W��ԶiU��8&�z��PW��9=�:�Ț�u�}sȸ�"rR!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��0
^�߽(�&����e�Y��R��go�'�( �~��U8L������n�� ηisȸ�"rR!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����q�<r�x,r��[�f�:&&e&���tP��"�h�j-���	�"a���7@"78X�˞�DG!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3wF�j�;�")$���/��Q!������sS�W�%�&� a�w*�{f�cI�yn��3<'���l�p�m~|��Lf��s)L��mU�����r��Ψ��F$��O�&�錤Ki�:�&x�.R�M6|��Q�՚�<����� f�+���c�����eי�ӿ��I�t~���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3K �n�^�b���?��/��'�fj��E�?Y��B��­��*G�Z�jvL�տ�זfEm	dmvPta!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3usA_�eP�2[Ӈ:t�y��ż�&/�� �g{��TV�yЅ�e�������g��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3"�(��t-�^/�?�\S/Av÷�������9�a'�!��)�Y*�&���1r��g��-,G�7�mEi$���0w����R�A�לA��P��粚������wb�S��V��\����Q��*�fjZ��9A
����u'���B��h���"�h7�o�/_�}v��؄aX܇5����`K<�{��E��81�� ����E����F�l����4v�7�ZSG3#z���=���M�>�P� ĵ�&�;G�7�mEi$���0w����R�A�לv���h���������wb�S��V��\����Q��*�fjZ��9A
����u'���B��h���"�h7�o�/_�}v��؄aX܇5����`K<�{��E����ʰi�B��E����F�l����4v�7�ZSG3#z���=���M�>�P� ĵ�&�;G�7�mEi$���0w����R�A�ל!�/�J�ٲ�������wb�S��V��\����Q��*�fjZ��9A
����u'���B��h���"�h7�o�/_�}v��؄aX܇5����`K��Oڭ���Ё��V+�
�c�~e͉�Xk����0���$v����_�'���qks�b��R���^.Z6�xI�7�а��"P�y�"'��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����P\�Ǿdj
>����p}�6�`s�$5׷!�Y@���v/�5��Vչb� ��o!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3BSyw1ߤ��,F��Ax�Zμ�2H���_���lV�v�bm�������8X�˞�DG!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��<�3D���iC\��"� vD��!���F�Xwux/.7��k'�w�����Ɔ�9$��i�m�����ܜj>��i6�0w�mo(���3�К��$B��Q{�C�Ɗ\CT20%�X�`<�`ۯn����T��%�B��ׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3uV^�HK9�g%�~�0ѝ�9��&�>���f�&�v4ȪP���W5�����Fz�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3 �y�NLAY>�>�w�I����,�1�%��;K�Jjףб����z�|�J��vsȸ�"rR!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��jy4��
����u'���B��h���"�h7�o�/_�}���2�O