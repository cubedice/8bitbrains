��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR�� ��������M7\F���r����&$9g8�M>PFWD#�z":���ӳ��_}��0w�\��8׋�������N���?��m��+�ڔ�wV��?��N��j$.:&R�nU���T���딣0&_���X0���2|	p��rw@	@us���)�]&��_	��u|��yq�`݊�|���"rG�
���}�\�bJ(9�{��r�H�����طǪ�`DY��YH\��!���1R�_ߥ�]��4�:j�l�,9��Տ�TG��1 T�V	�tL��	�<�A�}QP`��dpfVpb��#`^���w`qԗ�-�l��ǫR��p�� B]�pE(���B��|�(����5�%���(�-X�Ç�e�L|�w.j��6��H4�
� �AH��Wz�2���0Q����U~��{S�#�(9u��~�MUs ߼
�d��*Wq)e;�W_)O�l�I�"]�δ�� sfx�g H���'u��w)�SU��T�d��_�:�2�ٶ"n��v���uWTJ�Й�m�BM�Ɋ�p��"�U��b!��u�>o·,��8D"�s�z:�Ebzi`Ht����	x]�Ħ1��&��k���p�Z���Ǽ�5i�ĞX7�F@�4%���*ң3E���Xb޷j���zA&�\;��Ńi�[��1	��������k�8���҆�|n��l5����9�\���;j[���Yi��o?�M��;]��T��t��@�Lo���,,?���cu� �!+�ُ	Y��NL=�m�!=�y����h�}��(�'R����)*-1K�c��^�W�u���;�_Š;�������p<�������,�\gE�y�7�	����o:˨������|2��I�?5���q�xD�i�Kf���o�i��RL�a)Y/̹��~篟|����T�	ءc]"t�39����E�k8�Jlk�#�(�\��wŷ�8�2o��RL�a)��ô��o�~篟|��^��}�B���e�8�:r&@�G	���su�]bu̎��蚛y���\�4�s��)�]�.�Щ���qJG����A�LR����D��B��z�F��'�`�����G�Xp�m�!=�y����h�}�
"�k�'�2�;Y���<vF0���u���;�}����x)��>C7�`�����6���,���>]��|��ց��6 �ǽ�O9*]'U���k��
H���ܫo��RL�a)#�%Jd���~篟|��j�s����J>�C|��8�:r&@��|�)n풞�J��Jo3���_�z�^I�=�C����~��3>�I�z c��(�U����	x]��²9h����q+-���W��r�����G��F@�4%���IR.ux'V�vЊ�[-�T�g����g��5F��9��5l3߼
�d>ʟ;��BG-���K���RL�a)zAY����-�~篟|���"�9R������w�8�:r&@����:8E�#}�{��Um���P�����-�aeU��y�bK�D�L�	���RL�a)�ϕF���9�~篟|��=%����`O��{�8�:r&@,$h���o8�8��vD O�Y 7L��3K�<�#t����n��u�T�QU���2�B�~\$#����5[ |���>�
� �AH�|D3�MZk ��U�׏�.��GFUR�.�;�~�MUs ��\�j�ߩ&v��,Ҥ�P�X��AL��U;j~��`�{�y�ҭ��=�kM4v/:�
��$����aA�O�l/LC�awM��\�4�sg�oXx��UZk ��U�m�FƔXV�:Ѫ�2��~�MUs 7�_���4�l������RRK�*�C�r�O��C��0���M�<lbtsظ=��b@T*&L�5&#�u���;�;N��;�Dn�m��d�7�M�	Y֎�̖˄��O;Y����Gw��#�����]���Қʇ8[�r	}�n���M���E���k�8���҆�|n��I�� �r �/�tA(m~)i�d_�J�Й�m�X�LGA����w�F΁������m[�6��l�
��E�A ǢC���s♏��"� c��(�U����	x]�fX�eϝ(�Ua.{z_^��ҭF��8O �L#KX����/����}=��?�fO�ɪ
� �AH�W���,H�Կ+�H5H�*�k�-u�A�F@�4%������Ą���V����*�~�n_����uS ��������&�mN c��(�U����	x]�<���eo�l$�+���� �����Oh5Edɲ�<aED�2�Q�@�Y5M�e�o"�z�C�/7�o�H���7Ә��@Ő��tt=�L��r�O��C��0���df��SA`�/T-B�}8���u���;�'�� +�ۛ���p<�������,�\�H���UDcKE#�4*��1���l�,=�2\��c�鿷ŷ�z����~��M�{�ڌ�2¾'�UB�m}����������uS �����t=�L��^E�h/�����a畹�{�ڌ�2���-���t�VK4��i�;�t�!�k]�r�r����SU8��RL�a)3���ʉ�N	:.���nh��,+"<X��1� =��7C��H��;<��j6����V����k�FS�CO�����U���oG�gf��#u��w)�S��X3����~篟|�
�����2���Z��`8�:r&@��|�)n�bI�#�t�(HrdpSAHF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������V�e��Z){RQg8�]|�w�����N3|�}O���i��9�sT%lo�i��I�TY��"���u���KWʍ�I���~~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3ts�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S�7���I���}����E���ƪ�(����D�I�?g�fY�~�a���+�Uz�QL<(�P[H�������'SR����.�}|��ι%9T��7����+�Uz�QL�W*g;X~09h�i��I�?g�f�$��P�xZq��t�1�:�Ω��
�/�r}|��ι%9٤�2[51gyB-j&?��2�C�b��}Y���%�5�1�:�Ω��
�/�r}|��ι%9��oGo�Z�J��ݪ���AOge��e�IC�_�\�����@J
A��w|�<��y�~/r�I��
����&�ɬ� VU+I���ť1k�`��'p�@�I�?g�f��m����bi�ī*��I���0�1}Kط��4q������ |��J����>�Rh�XI։9x z�Jm]A�/����<.+6J!�p�ϵ�DE�U���!�`�(i3�b9���?̅4	������\{F˯�+)ƍ���� ���3�ҺIÙ=�H<z,Ҽ&�כ��p܏�<
DN�!�`�(i3JHn��z�_c)���8w�n���R�^Ƒ��!�`�(i3 ���3�ҺIÙ=�H�ς.fOoI�J��#Kl�Y�7#�xI��]n��JHn��z���G7���M{nnmCw��m��3��p���H����[7�d|���XP����@PVڵ��#���F�O��86�E����F�'n�^0o`�U+�PA�p�ϵ�DEG�p�P��g����=�b9����4�6�t�8֩]=$�����k!��V�_g� ���3�ҺIÙ=�HF���m¡fÁ��/�6�_�"�,�>E����\�v��_�R�G��W�$�qx����Ѱ0|]<w:�,ԯ���gn�J����� ι��QG�����U��!�`�(i3зq8�Ј)w�<�_N���i�����Y�V&��A��.D0I� X�1�зq8�Ј)w�<�_N���i�����Y�V�~G���7ht��}jзq8�Ј)w�<�_N��}��|�d!K-2�E���M����A�m�(�� nU�IÙ=�HF���m¡vuƇgv���6�=]A��O�T=�4e=��-��̰S����T<؛L�kT�䖙�Dys�зq8�Ј)w�<�_N��k�����\��>O�S�e�}�	��%�Y)���N�No��c��u�zL͊�q���\��;�,�����w�=5[������#s{��'�-r��|ڑ�H���o���&�t.�}w�n����|��T�5�d�,W�� nU�IÙ=�H��'�PD����
q<O�n����9��#�B�sYC��\�v��_�R�G"����?e��G�K$x/��&��닞��D	��U�l>o��|��'�njVfV����x�%�$����{v��G�K$x/��&��닞��D	��U�l>o��|��'�njVfV�*lZ����]V�H7'�5�}�]���!�`�(i3=]A��O�T=�4e=��-f[� ��³��w�[��C��!�`�(i3зq8�Ј)w�<�_N �VL�(\F�c���$/���i� � �	{����0�&�ͭ"�,�>E����-��%Mό���.��_F�k-�!�`�(i3c��Et��q���U��;���)"����}�����|g�Y�'���Xw�,bxqX��9��no��b�:/z��]���c�A�L'G~��6�7*���T��
����ѳ�T�\ �͘�f��p�b�z'hۉ)��d�7�q����B['u�E����F7G#+��\w��0]�r���h�0"�,�>E���TD��ό���.�q�\E��0M7$���c��Et�Y�{'%s��.|Z���I7��-5��6��	���`y����ꢤ�Og�[N�&ѐ�����
L'���Xw�j�7��U����z~��6��	���`y����*#�m z����Z��o�����
L'���Xw�j�7���=�$�ЭU����z~��6��	�\�HP@�a%=dϖ�i�@O�x�7���q�©��L�=ɐ<c����4�Q��ņD^�NË�����8��z{��E�EYZ/�矘��-n��I�?g�f��m����bi�ī*��I���0�&v��p:ڃ���開Ŗ6$\Kʯ!��}Y����
_#@��#	T�d����'3ˁ�ֵ�r7����ݸb����b�N��q��p~E�>@	L���M��fk^,��rk��4�o�r����_��A"�U���w�c*����_|1&�����'3pk~������8n��.V��8�nT��8&���I���8|�p�ق�4?}�\�����Ք�)�"1tSjv���=�gw�⽒�#9NS��1	�q��p��'1�F�NQ?M8�f2o|���P��4Q��@���ݚ�Н��x���	R����>�R���mK�g+Wx�Ա�%��ݚ�Н������VVw�⽒�}�\�������9��
����	�|��!�`�(i3�<�I��y�G��C�m��U�E����&��&o��ǈ�A0
���5Q��!�`�(i3�?�JY�)�s�[7��!�`�(i3)�{6�U��$f��_Ub�F�S�1 ��?�JY�)�Y`��jD4}�	76�&��A0ok�����a�"�_���3�<`c������偋:�Q	Q��|��=+�	QH�&{�H�u��m9����L-R���KO����1@n���Js}����R8!��vp�P}��O��ꅽ52����$�Qu�&�<��G�JHn��z����_�K�}��K�&`ZPյ[+8��x���	R����>�R���mK�g+Wx�Ա�%��|#HK���\r([.<J�M����!�`�(i3�R'cf�� ��B��h�W. �9�����Yk����Aڬ&W��K��1?�j�EH�RtV�^�y��j��k����ï!�w(�y?
�:qEp�;�P�t�5
�:qEpCt�w#��@�����fĉ>99��A0ok����jVѭ@Ƹv��*Qx���x��@�2N����RUS�f�:䩒=]'ʥ�nr]�b�N��r�t�L^��޿���Y߼
�d\?�����k�O�%�d+�����蠿����d�Uf�揆0�б�d=��¾ȼ�}�٢�% :�ǒ���K����������a�"V���9س�"�<��E������sc�v	I�����F��O�C8 ����C�ӼGt8��Pip<ɯ�nv��2������開���Y����Ů�;	�nw(��=����$?���*{ٝ�,���8! ,��e�ŷ֗�e�a�i���S=GϦ-�:QT��3��L���*ތ�@���[�Bf�^:.���us�b��v�\��JHn��z���!>����8���ao ��M��_(����@҄���G��A"�U���w�c*��t+��I���XP���ʥ�n2`qd�#��Ӏ�`,9�H�WMl༗g##���O3?ӽP�y�[��(��Ƹv��*QxR��9�H�@͗��3��}�	76�&�R�V�"�0ɶ37y�����:������	���Nt0���l���r�z�dQ���߼
�d*��+��u�׫A|O����/;^��(@v���N�l:�Brq1��B�ce����:��'��Q�f�G\&��g����開&ޗ����^��/�/m�d�ů��z��_#Ԡ�g��2у�ӣ��[���b9���M��A���"�g��bc��[�Bf�^:/��T�n*�N}�m��{B���T�D�}�+�r1D��y�^��6�Rsb�d"L�%K��ͪM$յ[+8��i7N�_�Ar��� �nק���!�h]��y�Q?M8�f2��֖+�)�#U#��F:җ�S��dZ#'��� h�ҩθ<�I��y�f7$=�0*՝� s�#���k$ Uc��͘���sjl̓y΢�Lb&X��0d�4� h�ҩ�֭�h��O7�aO#h���}Dq�f������!�`�(i3T�zU�k���n��u��r��!�`�(i3�zk���~�-��:��o�R����8N�������aR�!�`�(i3�����!�`�(i3�<�I��y�G��C�mđ�e�a�u�!�`�(i3���F��O��ݚ�Н����F��O�!�`�(i3�;b�-�2��;�P�t�5���W0�]��x@�������a�"�_���3� �n���.�c����Pw�������#p��H��R��Y��(��v�r��6���֓�Ӛ}���9I��@��p�m~|����j(�F�H#
ZM��,Gk����1�~��)�K�e��T���u�I���bU�򍬓BS���U��*ң3E��_(����@҄���G��A"�U���w�c*��t+��I���XP���0��QM�Dx�ܰ���開���?�`�7Ue�B ���
��]k�y�"�V��5M��z�o$�S�in���),��9��"!<n��8��dט�w�����T�ɑk��!a�tc�&ck���������IÙ=�H�R�����|c_�m��ġ��,;�ŝ_�fu��w�K�	�<���BSG�p�P�Jٯ�n
�5����`K��M���-g?���ų!�`�(i3�b9����2�u|�*�7`����\Z��K���\,��#t�z`0yM��^��q�3i�<�-�p-ʅTV�����$��Xo��yذ��t�H�MPq6.!�`�(i3%Ah�%4
>��XP���ct�:��RE��W� y�T�v��1���2���I��'��q�2�_:��p\I��� !�`�(i3A( ����_�h3��{I��Z��H1�$ԠI�*U2��53���>G�T!�E����F�'n�^0o�VU&ZM��9��"!<n��8��$��Xo��GR��)�hvl��9�h �=�%Ah�%4
>��XP����&ތ1*[,�v���P�V��>'�o��&L���W=D��'n�^0o`�U+�PA�5����`K'{}yw~�귈nIg�R���]6���b9���P9b���dט�w����4��}>0�1ۍ�h �=� ���3�ҺIÙ=�H������/=3\H�d&�.�_�L[� �h���Z�j-J���\�v�X�zgq��p�m~|��wʞ،:쉎���AK}�p~z�r,Ln��S�W0�T��:*�����
	�7F���I@1���t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s��.|Z���I7��-5��6��	���`y�����g�,P�n�Ͱ��Le�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cUL3�X�j�>&�&i�"j���b7���Øf�$��Xo�U)+N��e�J�Pn\�=�����JHn��z�F�x�aK�k��Y��)ё�H�a)��dט�w���f�ܗ��DX<�c>1K �:;k�+��b9����|i��I��yN��7��aq��hx��t�#���Fν��E�p�m~|��;~7����WF�r�f�t a
��Vx^��\�v��\aьIR=���|�F֣z>Q�Q�<%�a����D�K���g�,P�n�R<�����\���^�W+`�x�oP��@t�&�e�5
�`#_G�쵄����T�=�;^�6#9���k��$a(􆿳�ټ*w2�56�5����`K��M���R'),��`�?2{���zL͊�q��*
�DWo$�}��M�+�C
2����Ol���$��Xo�e_�d
���ݪ��1#��Z�����XP��ȗd�uY��K��T��p�AqeGfB����N�e�8�ʫ��;ƹ��:i7s�9���o��S8���/=u	Mk��!a�tc�&ck��*h���'�a�?� Zh�R?�R��n��am�Za(􆿳���2����.���N�e�8�ʫ��6���7s�9���o��S8���/=u	Mk��!a�tc�&ck��*h���'�a�?� Zh�R?�R��n��am�Za(􆿳���2����.���Nihc�ؓ;)�;ƹ��:i7s�9���o��S8���/=u	Mk��!a�tc�&ck��*h���'�a�?� Zh�R?�R��n��am�Za(􆿳���2����.���Nihc�ؓ;)�6���7s�9���o��S8���/=u	Mk��!a�tc�&ck��*h���'�a�?� Zh�R?�R��n��am�Za(􆿳���2����.���Nihc�ؓ;)Ve��˅�O�=�ͦ��r)��ׁ�a\Y����+���LQ�g��U-�e,%�0g�������DzL�����A@!�`�(i3��?��(��I@1�ؠ&���Z02��`�z��Y��)�D�YG�9���,D�K��D��`'Vp��U��E����F��
��D&e�2l��4��a��se�ξ���I��RhF��?�1�{}�
�?�&�z���@h��,��!iJ�p8�(�E;*�}Ւ�~ܔp�l
d�R�.��On��M����A�m�(�Jٯ�n
�
�CӞD�+5�4��c�M�����U,�(�)8⋌�U2ރ�8���/����,D��8^a�F~��^x��G��ʡ3��jgZ鎬�������(�����y>'MM귈nIg�R݃��x���g��U-�e,%�0g��սÕB\�6NYlԘ=�!�`�(i3��?��(��I@1�ؠ&���Z02��`�z?�R��n�#ٷ�Ef߸@����gG���:���U���;�'���Xw�j�7��g�]@n_���?3MN�-���8���/�I����"�]�N��&�|��sQ�G�O+�|��p �>�Y�{'%s���F���-�'��0�=<MW�-}�	mp,��_А#�<om��Pk-� �!��.ᬵy�����u�4�����p���yN��7��aq��G�n���t�;���NK�E�l�b��ƍ��o���Øf}�
�?��Y�Y`$�E�.1p�Y,_�S�
ut�q���U��@����gGz�I�`�M�&�^���зq8�Ј'���Xw�%G��ly����DzL��T�B�X
ŝ�2(4`�'���Xw�j�7���ļަ��P�of$��D�_�k�W�A�&hH\�T�\ ������q�f@x9���7�7s�9���o>��l%i�-�n~�x���p�	O$�]�!��8�$LQ������N��H���9����}�ڍ�xZ��j�
�&�j��1�a-���7a
��r��Q��Y����2����.���N��H���9����҉}%xZ��j�
�&�j��1�a-���7a
��r��L;Л��|#9���b!��u�j2�K����S�p�ɒ�[��&�j��1�a-���7a
��r��Q��Y��ټ*w2�56ݓ��E�/�������� �mDL�>��0��Q]� _m�jp=�>��o�
�v�ξ���e�J�Pn\���p_U
#i;��#��F�r�f�t���ӯIJ ��`y����@����gG�DI߃���iA'R�	md���{��E����F�R<����z���踫g(�r�x�y�Zgl�k�����դL� s�j8��L���N���"�L�6yd(!�`�(i37s�9���on�-�6��
�jW��D���M���o�G�m�?�5:�7�+pVx�%L��W��_�ړ8���/����,DTc�~y��i���n���g!�`�(i3"�,�>E��[��Q�՝�i�(�S��]Q�I����踫g(�r�x�y�Zgl-�g����,DTc�~y��i�����-VL!�`�(i3"�,�>E��P"G�wk�P#7!smWF�r�f�t���ӯIJ ��`y����@����gG�DI߃����t��!�`�(i3�E����FZ鎬�������(����S� ?�0��E|�,°������R�wX��}�
�?�N��	�Ȓ�cЉ�M�C9*�¢���lJ��튝�b�Bϱ��R<�����á�~O��L;Л��|#9���b!��u��Ɔ ���.�&�?��¡J���a߲��+�J��Y�{'%s�h�v��[�x�X���+���LQ���"X��[��Q[R�7�B'�P���h��LwN����ڕ���V�6IWJE�r���秹�3I^�v�%j���x�;��ԁ[�x�X���+���LQ���"X��[��Q[R�7ݓ��E�/�����sc�̆�!YV����-�~8;��Ҙh��LwN��j8�U� %G)�Х'���;���N� �vf&}�
�?�N��	�Ȓ{A�dha#4����ʴ5��ǳ%Y�杌b�Bϱ��R<�����á�~O��L;Л��|#9���b!��u��Ɔ �����O�����C�1�r5��(әxZ��j�
�����1��;-;*�7��;mQ��8���/�H/�B���L���N�b�'Beͧ��&�~Ly�1O�r^Л[�l\���$����b�m��,���b�U�J޿�ġ��,)@����Sb!��u፵mp"�o��}��u@:��/y��g�'b�t	�U���C��O]r�<Uee���nH�W�]��fM?R�^Ƒ����"X��[��Q[R�7�
�CӞD��~VHx��_��x�7s�9���on�-�6��
�jW��D���M���}a�/�kj��NI�:7�N�5�%]���a(􆿳�p�Q��j_YK�}_�zc�bK�s�} Oag����W{~�85Zt���%�]�
ƇBHx\�'���Xw s4S�'�i��`�z������1:#�j^�y]/�qF���ӯIJ ��`y�����g�,P�n�BL�Jx��e�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cUL�f����Y>1�Z���=��L;Л��|#9���b!��u���t�f�2E���n���g4K�)s"���݇�T%{�;���E&�0�3uH�,�7�%�a�A�m�(��X����[�ǈ���?5���q��6��v��o�>P�2-i_��]�v*&��A�YHm��G�m���+k&v�IzZ鎬����
C��8q��f�kN�ı���}J�|���|����S���m|�U����z~���ӯIJ ��`y�����g�,P�n�i�_:�ܷ��	N^�U��J��"ї>п�p=	�˳͠m�xW��9u$d9�cx�S�����S8�����NlU����z~���ӯIJ ��`y����@����gG�Be|���������v)o21��I�L&R�B���B��㎏qló�{��]z�����Dɵ�p�AJ�e�$TA�𼀅@����N��"��=���b>0���`!�5����`K��mV�T�D���ɻ�������� ����U�P���4��=Z�˂�hF���H#
ZM��L~΄gO�3����?��.�����<	: ���@89��i���"<璋���n�4�{lGD�V�Bf�Nd+l�Yҽ֗�2�0]�J�$��Xo��LL}�և��6t�.�!�`�(i3l0��F��jY_���P[!�`�(i3!�`�(i3�;C@������M����A�m�(��`PV��yN��7��aq��hx��t�#���Fν��E�p�m~|����
���լC�r�X&d�X0��ތ�@���[�Bf�^:{lGD�V�B�}q4!QA�Y�x΁�)�<u��R��0�z}�Jv��m��}�8P��1prB%�?��Z�z�c([p�m~|����
����~���e�)qP@L0��Uތ�@���[�Bf�^:{lGD�V�B�}q4!QA�Y�x΁�)�&ޗ����NW����#�ٝ�z*�[��5�-Q��yN��7��aq��G�n���t�;���N���ke�zEp�m~|�����Ҏ|�~@�\��!�`�(i3�d�ů��z��_#Ԡ��@d��שI4��欱���j����w��G�Ŗ6$\Kʯ!��}Y�,����f�� l�o�bw�g���pǓ#5����m��3��p���H����Q#�?���;���N%�:+W�5����`K%{.�V#?p�&���A�=�א=ͼ�\�v�!�`�(i3!�`�(i3!�`�(i3!�`�(i32���s���(���B���{�T��Õz����o�8�v��(f�Nd+l�Yҽ֗���Z��*��w�>��p�&���A����0��V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s�O��W��W���}���i�����dq�8���/����RY��Ɛ�<["���܁�_�4�|�D�{�W+`�x�oP��@t�&�e�5
�`#_G��j�i�+-ڎ�>E�%��*d��:=�;o����׋��`y�����g�,P�nv�@[�JJ�-t�A�ݔnb��M\A}����gE������e��m��3��p���H����Q#�?���;���N��'?X��vcx�S�����S8�u�?�f�Rv�@[�JJ1��P�M���L;Л��|#9�����:�<�L�E��w*e�΢���vD�:�d���u�hF�
��ӧ0�=<MW�-}�	mp@�s�p���.ᬵy��k�t��8*l�J;�R^kAO��t��y	����F��،°������R�wX��KM���d��7Syv�J�Յ!��4�$��O�&��;�L���9�D_�3���U_�+X�P��y7Syv�J�Յ!��4���_GI�� bL}b����*���G��h[74�[U�9�V�6IWJE�r���秹�3I^�v&���xzvL�E��w*e�΢���v�R�U�S�cb!��u�d��}U؄�k]m��!�`�(i3GYs��$;��H��,x,����ar�<Uee�N�����H�OM��`�@����gG�x���يj}c��ko#�D�d��k��X�o�!���	����}q?H^��2踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��{�j��<�ao���wE���Ov@)�l��0�L�E��w*$��O�&���f�kN�ı*�7`����\Z��K��tH۷�ݫ�/h�5�G�Gd��}U؄�k]m���yS&E��1GYs��$;���$���M�;�E,0�ΩyO^~��M����A�m�([}�@��L}�
�?�v���,Ͽ�2[QvA�ͧ��&�~Lb�W�[*���G��h[74x,����ar�<Uee�N�����H�OM��`�@����gG�x���يj[��m�UZ���,���X�o�!���	����}q?H^��2踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��{�j��+�g�>U�6���@)�l��0�L�E��w*$��O�&���f�kN�ı*�7`����\Z��K��4����/��.������FD>�v��t�損t�5�v�@[�JJ혮��ר{lGD�V�Bf�Nd+l�Yҽ֗�2�0]�J}�
�?�u����p�5�"��[�BȒ�0^M�b�W�[*���G��h[74���E���:��`�z��Y��),�B۸��L� s�j8�-D���6	���� �[e�~' Y�]�7Syv�J�Յ!��4�e�p�������
��M����A�m�([}�@��L}�
�?�u����p��8��V\�J#�	g��b�W�[r��-�W.��@��i�=�f�kN�ı*�7`����\Z��K��4����/��+w�7�~�Y���Wql���B	�A���v�@[�JJ혮��ר�bl�_�p�ξ���I��RhF���k��76����,D�ʥ��G�M��KJ#�	g��U�î�D�p�&���A��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u�zk����G7```+��֞8�V��GYs��$;��H��,���E���:��`�z��Y��),�B۸��L� s�j8�-D���(���!G�{%(Zr*���P�e�b'���Xw�"O=��踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��S�8w?�s^��ɷ��e�ݲ��+�J��Y�{'%s���gt�͓�ξ���I��RhF���k��76����,D�ʥ��G����9�~��� ����=�^�)赙 ����/?(��=՜r�<Uee�N�����H�OM��`�@����gG"�t�'ێ��0+��?l�/��X��n`5�fK�gh1�͖5�Zz2|��M����A�m�([}�@��L}�
�?�Z�,��#�2
��e���.��;�#*�u��6�gh1�͖5�Zz2|��M����A�m�([}�@��L}�
�?�Z�,��#�2
��e���.��;�#]����),Y�{'%s���gt�͓�ξ���I��RhF���k��76����,D\X��!��x�D�Re�@oX��U�î�D�p�&���A��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u�o� c �R�%1���%�㴭+�JGYs��$;��H��,���E���:��`�z��Y��),�B۸��L� s�j8��h��)ew���m��@oX�� Y�]�7Syv�J�Բ������sl����?r�<Uee�N�����H�OM��`�@����gGچ�����F�f�J�㴭+�J��X�o�!���	����}M�l8�	
ڶ�@d��שI4��欱���j���-+��B�G3�+��m\n�v�ĺ�֦�w�#d�7��h��;	Ɛ�<["���܁�_�jZ"]�Vp踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀŻw�sH,@��@R�^a���<�"@)�l��0�L�E��w*e�p�������
��M����A�m�([}�@��L�@����gG�x���يj}c��ko#B���T�Luv�@[�JJ혮��ר�bl�_�p�ξ���I��RhF���k��76����,D�x�/��Y#ѥh��k�~ҤƐ�<["���܁�_�jZ"]�Vp踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��{�j��<�ao��<�_@X��GYs��$;��H��,���E���:��`�z��Y��),�B۸��L� s�j8&��f;�P䒡�3���α� �m�Ejb�W�[r��-�W.��@��i�=�f�kN�ı*�7`����\Z��K���^���?���)�`E5kUx���6Z.��0�W'���Xw�j�7���R<�����á�~O��L;Л��|#9���b!��u�fePh�����=�׸��d�٣��c�A�L'G~��6�7;-;*�7��;mQ��8���/����,D�;����;��|�D����Q]� _�rs�i��@�N3,(�;^�6#9���k��$a(􆿳���2����.�N��+�j����tL�f��d(s��d�٣��c�A�L'G~��6�7;-;*�7��;mQ��8���/�����s�c�����gv,��u(q����hc� ��;����Q	2�1����޳va�{����PD}#��ů��èV��֖+�)�#U#��F�E�P"��Wx�Ա�%������a�"��w�K�~Ҹ�`*N�ǁ�f�T���j�ʾ+)P�c1�(����C4'n��=?���͞��>(�J5����@|������]��R���}��M�+��l~�U�{}��*�}�	76�&�� Ӗ�tJ��K�]���!E�.tik&�#�P4ǲ ���"��|���it	�Tߦ^Cg��) ���3�ҺIÙ=�H槑��gL��dn��A����QߡN���ޛ#F f�Nd+l�Yҽ֗��$��'!�߼
�dV�I~!���(����C3��o��=�1+�AK3G�4W��(�!�>��y�P}��O��ꅽ52�����8-|�D<���K<�%�/��Z>L�<��˓��>�X6�j~ʮU:�W����vcy�3�"��+W���F�^��NP!��"� +}Z�"��%o�N(��~ӧ�1�Z���=�Ζ�,�Z{ �=�%�*�]�1���Ě���aT��3G�E��ч¼xE���8�|`��P���(h�(�
�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����sC���"��|���it	�TU����z~+Yi=��o�IÙ=�H槑��gL��dn��ATN��,��n��i])<}�
�?����*�t��v+�/;�d�٣��c�A�L'��Gr_���GF��a�1�Z���=��L;Л�����Øf�$��Xo����BɊ�y�+���LQ� ���3�ҺIÙ=�H�z~~�Y_" �g8Yw�
��vK���w�K�̄�Bq���ZLN�	�� ��˽��r�Q�gL#A=��a��'�-�O�Y�I�4];ˍH��KD:�}��0nk��ކء�Ch�1Ǥ �)�?�0��Y��W���U�dP_\G�7^2$S�6���f�_)fxg��pH���0�Ҋ@)�t�d�f�rЄzɳ�B��,��C-2�^���ij�IROgn�t���c�&�<�o��H�,>��*�:��I�}L������@���t����N@<����fRD�}a�/^�yQA��D,��f�x��r�@����gG<F��̎ÆWw3i�|�зq8�Ј'���Xw�j�7��Q�%�+2�ƃ
ᾆ�x�T�\ ��i3�|)sՀ@�g}��c��lmR�S{}"�,�>E���]�!����w�Հ�	:ү0CAe[u�;0�!�`�(i3�d�٣��v_���Zo�����n9�c�!{p857s�9���o��S8�/ #O�)R�^Ƒ����"X��[��Q[R�7����n9�jsrCm�k7s�9���o��S8��Ѽm����wk����\����|ݔ�3�(n�'�PW���[f���Øf}�
�?��YN
��)eS���c,P"G�wk�١��	;q�J�� m�h�5,Wlr�r%)cA�z���a�R�wX��}�
�?��YN
��)e��g.��P"G�wk�١��	;q�J�� m�h�5,Wlr�r%)cA�z���a�R�wX��}�
�?��T�n��a�S���c,P"G�wk�١��	;q�ew�:��w�<om��F`���G���`y����@����gG�;�m�PV|�LOo�xZ��j�
�iB{�Z�_�+��tI�F�;���Nk��}�y:�8���/����,DJΌ�#<�F��6�q��T�ٮ|�,
���1��e0����yN��7��aq���E���ss�T�\ ��i3�|)sՀ/��{��`VTҝD!u�U,�(�)8���0y�	�l�f<Rqا �GR��shbvk~�#xTU]O�d��g��U-�e,%�0g���g���gQ��9mh��n.�G��J��\[$Q��
�̞��>��L�溥����v�8:�x�3�Aga(􆿳���2����.�t������H_��#���1��_*|AԢ�a\��F�dHB�Fvͧ"�f���-A�¤�x.�Knq�z���a�Г�����]���3;�7���c�	4��t�f�d�٣���N N�S�qg2�K?\�2�q��n`5�fK�\w��0]b!��u�#� �,Wɒ��r����q���U��@����gGNc�&�Ia���`M��
Z鎬�������(���j~�]�������:�.�& 5f��e�T�\ ������q�f@b02�O#h�\�̐�]�!����w�Հ�[�=�5x�����P"G�wk�ED��G��|#9���߼
�d�Ȯ�\	b1X�7�o����I��8�M�$�愉V�Sup�xg쬉� }���n4s1��7�癆cg3bQ=�3�� �֤D�A�f�8
��u��r��R�@�6�֐��s�;�9�����:�.�o�J��h�׮	��48ܼ�P���#�紩$�_�B&��p�)Y����2����0/ܤ�(g��V��T�� v�0�=<MW�-}�	mp����"���;���Nå�a1��Y~�y������7��[�G���P��w�T:~�f��ƈ�<om����[��l_1���~�37y����~#f���-�o%��5��/dV���(��g.Cf����)Y����2��ļަ��P�5��/dV�z~~�Y_"R�W�uy�cs;H��yN��7��aq��͹��e�[�.ᬵy��H0@&ɡ��Օ��qvdЧ^{�j�E�i�m}6O�D mWN�&�ҙ��Cm�-H�h�Usdx�������aR��$��Xo��4�!`��] �v"�O���-�SIÙ=�HQ}Sٔ&Fƒvof��l _TЬI�]���3η�H��:�-).^QQe���b�!�`�(i3q��T�ٮ|�,
���h���J	�0�ȷS�J����Xa(􆿳���2����.qg2�K?\���a{�5���u�L�!�`�(i3ғ�vq�\[$Q��
�̞��>�nQ�rV�}!�@�?0a(􆿳���2����.�E ����$,K�9+�/���p��8�{�����x z�Jm]�#�;� �@����gGP���Ʃ8/Tu�����_&��������]�!����w�Հ�JX-�ܶ�0l�x����b�'Be��
����ѥ"�8���q���U��@����gGP���Ʃ8/Tu�����_&����=/����67s�9���o>��l%i�-�n~�x��Nh���W<˥�'ܤ",^� ��B���+�J��Y�{'%s�
>���d&�.�_�L[� �h��MN�-���8���/����,D�8���Q׆��p0�Ĝ(�IyI)wf�U݋s�n`5�fK��0z�cULA6{'8�0��9gP�U,�2������}�{q-Tjo�R�wX��}�
�?�&aD�4�X�X�>c�.A��I�JZ�d�٣��c�A�L'����8?�o[L��h �=�.�v�L#�?��Q[R�7�n~�x��Nh���W<˥�'ܤ",�X�G[�!�`�(i3�n`5�fK�gh1�͖5�Zz2|��M����A�m�([}�@��L}�
�?�&aD�4�X�X�[RP� .���j�#-����E����FZ鎬�������j}�c��`�z��Y��),�B۸��L� s�j8JX-�ܶ�0l�x���
��e���F7�GhzigzA=v)�n`5�fK�gh1�͖5�Zz2|��M����A�m�([}�@��LJ�W��7/��)׺����\� C&����q��Z���2%�ɛ'���$� c%ij��d���0y�	�l�f<Rqا �GR��shbvk~�#x ��M��.ᬵy�����L7�oa(􆿳���2����.+w�7�@�Af8�ٕ��(�W�!Ċ&��/v�K7%'���+�J���q���U��@����gG���U�\ʭB��2�k1�h�H��*/v�K7%'!�`�(i3�d�٣��c�A�L'��$;-,�J�d�@q�2������}°������R�wX��}�
�?�u����p�����+X��FJ���-],��%s��u��at�kZP"G�wk�١��	;q}u6��\����m��3��p���H������7Pr��ġ��,���=�8���/����,D���S�D��_�W�.��;�#�E���_	!�`�(i37s�9���o>��l%i�-5�e`��9����dz����NR�p�+yG_��\�!�`�(i3зq8�Ј'���Xw�j�7������1H}�ɐ��/��HM���#ga(􆿳���2����.�>��왩�/Tu����W`GU�!i&G�\��u��6��+(c7s�9���o>��l%i�-�����bpA���3A�n�+�sQ}b`�����V@���gx2�n`5�fK��0z�cUL0x�?����z'/)�� 0�s]MN�-���8���/�i�V���kP�?��ԭ���|��q���� $�~����pk�,�Y��S��q������5*g]�H�X��%�N(��ڈ+w�7�@�Af8�ٕ��(�W�5���^�u��������+�J��Y�{'%s���gt�͓�ξ���I��RhF���k��76����,D���S�D��_�W�.��;�#��f��w��]�q�7s�9���o×��̙�F�9 }�m�f�Nd+l�Yҽ֗��i�ܰAb!��u�R��ak����`T�ҩ�	r^W	��s����a���2'���Xw�"O=��踫g(�r�N�ǁ�f�TpD��ZOUo�$Կm��!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vco ��Z�� ќh~-s/�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcj)�[N�|+_��'5��޸�~}	�U�&U����o����ϯv���&q��v~Azx�ǁ�j��C��][�j�r��e&�2��&����_`��ƥ�Z`���������B3$�#-��o� �Y��*6���SK���B��C����D�%ح�e!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}��V5VM�d�/|�;{$�WaU�����W�1� =�cw��혅vº�w�⽒���M����A�m�(�#W�U��ظ�d���!i�^Xe�����'HY-��Yk"1/s�\"�����p"π9�^N-~H	��`��,\ަ�It��+g[��v:ι�Y�0��E|�,VK�5��&q^�`
�c��><�$�"���$�(���B���Q��ǺΕR��ӟ-���N�����W���`moF˯�+)Ƌ��_��F˯�+)��&�C�/S��ك6
��^H��sp�]3t�ݚ�Н�EfVNN{s�ܱ?'�EfVNN!�H&y�i��[��C���������a����"�$,\ͨ܉p����O,8�ݚ�Н����D)���:��]]t}c��ko#��Uy�~��</Sn��'B�ɏ� ��U�Ͻv1a{J�v0�A��c[�л���7�Rz(��g��}#�U����5�W@�2��}���C�#�J�{�V5VM�d��m�.j	f�?ǉ�=�Aɀ��{��W�ł)w����ʮ��?G�+5�4��c��W������Ri��!�`�(i3k/�z�xEQ���*[UxG!�`�(i3�չ�Ad��vIn���Ԥ�8!7��%G|�<)���WR���jٵ��.ᬵy����*e@�__��s�֙7�}�!��e��E���&%�=:����c�/ROU��Y��),�B۸��f>x�:	�W+��W�s->m�9V��Vv��8>��
��
 %���'HY-��
�C�Ʌ��HW��ݚ�Н�R�7h�,b0V�u�Q�ݚ�Н�¥������]n��-��w¹��<d�,��L��!�`�(i3��.��֞�������i��D��;jQ�#���F�;�@"��ݚ�Н����8��T�h���}둮j\����C��rR#K�p�ݚ�Н��K�^��Q��G�S>\.�!::tm�0�i.�9!�`�(i3�2*Q=F���q/���<�����7
!�`�(i3�dv��oTN֢&@��&!�`�(i3k/�z�xEQ���*[UxG!�`�(i3��|��p��PIQ#�C,0�?���!�`�(i3��9��稕�a�/!O�f�?ǉ�=�2��}��CϾH�)�V5VM�d��m�.j	f�?ǉ�=�2��}���zgm##��V5VM�d6��0]�1�v�9�ʅ.�g3Z�Ǵݵ���pÓ�}<�ž_�F�Tq��A��s&?Z�l�(�u��@t�qP�V>tI��RhF����u�*��?�d���&��ݚ�Н��V5VM�d6��0]�1�g�)�I��#�r��8��ҥ�|HN��R��?�d���&�Tq��A��s&?Z�l�(�����0`;�V&S�b6j�"Hsކl9�p������l��Vj�Ra�m�,�*��'��ҙ����
�Z�S$J�	�LÆ�c�9ʼ��$l'>����J��:����9�{�Jj3�a�5@�i�QR�j4gM�+5�4��c�� D�_\HN��R��?�d���&�+r�^4Y�BM�e�x�U3u��� ;��|B�.y7bژIl���o���8�:�����zV���z%�/��Z>L�'��D(M&��w>��Y��$1&O� �k�3��6J�Ko��ih�|����
�Z�S$J�	�LÆ�c�9ʼ��$m#�P�J��:����P� d�c�.1p�Y,��J��ۍb�o��_�Rv�䩲$����tb�����+�^n=\f�5>����Db^�.1p�Y,0Y�X��f�\���F�`yx�>�+X�M?��y�!�`�(i3P���x�NS���U��[��c��3|v��Eb�z'hۉ)��d�7�q�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�s�Yls��8��GM��-����!�`�(i3P���x�NS���U��[��c��5H)�c�8Qł)w������U+��_����E�ł)w������U+��_ �2��9gUS����a$�/ϟ��7�4�.1p�Y,+
���Q�"���Urܰ#y���:5A��pfĉ>99��A0ok��fĉ>99��A0ok��W?�;�끓��~�Ly�$�|�m��Z�f�WM8}�	76�&�;��|B�mC�8	�XB�����C�����tP��b&�\JG8q.j<��IZ��x�,y�#���F�F��b�\��Se���7�}�!���V5VM�dC��6�g����5�ź�+���*#nC��6�g����5�źP�?v�l��+�ϸ�i���U_&�W\�a|��sQ�G�3��ݹ�w5���i�w�R���y>��yСQ=!�e���26}�i���:I�#��y�$�|�m��=�_�7V�o��_�Rv�䩲$��GQЌJ
��`���φ��<�6��ߙ�[�>	ol�~{�Ž\���F�`yx�>�+X�M?��y�!�`�(i3��6J�Ko�����P��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��y�!�`�(i3�<��7gҠ�(�2ʛ[�q�ܦ	&�P��k�Ӿ]ܦ	&�P��UB�I'9gUS����a$�/ϟ��7�4�.1p�Y,v�)�DZ�ϟ��7�4�.1p�Y,Q� R��F}v���۹�
�:qEp�;�P�t�5fĉ>99��A0ok�׹�����A�;�����[�F$�kj���6J�Ko���zX��-Z�+�ϸ�i$x���z*�7`����\Z��K��rt=ٝ��b&�\JG8�j(&
M�K�<�
�d�ξ���'�̗����
�t�c��5�O�%E#Pc�{��lq�<b*�_���t�T��?E-h��`f���s��6}���iI9�o«IX0F�M��6J�Ko��hm�ko@h�H����Qw�c4~Nr_�mS8<�n�ݚ�Н���� ff��X	n�ɺb_X�XV�b�z'hۉ)��d�7�q�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�s�Yls��8��GM�`�(�4�bł)w������U+��_����E�ł)w������U+��_ �2�Ъ��tj/�՚�-����!�`�(i3�<��7Nǌq�p�IC&��b��mf-W�c��ǳ��&�!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rG߸��S�Ȍ� �Q$j�sP��':�HN��R��?�d���&�x�����<����՜����� ff��pH�x��]'\gWg��	�Z�kfc?�#	*]]�iI9�o«IX0F�MG�k�P[�;�jmT�#bs��2[�a��o���H�RtV�^P���x�NSB���j%Ř�I4��欱���j��������my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�y�}�6f&r#o�]�ʄ�lZ#s��kgҠ�(�2j�y�`CrgҠ�(�2L���yF��G��Hb� h�ҩ�,��G��z#�r��8ߞQ���l�N�����K����F?Tq��A��ske��|ξ?�R��n�#ٷ�Ef��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;���z��O�Q��D��y�t����M~V��	��y��E��D�VvA#&��Q��r��`�@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�_L�oe��Em�Ԣ�+d%�4.P�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcN�H"����H��X�����k楊HaU$kX�M�ŗ\�'	�?��[n8�A�A���p������'HY-��Yk"1/|sL'���oֲ󄰊�������M�����%kR��������֢&@��&���o)�]r k�|6�8NU�:|������k!�M�Z���	f�?ǉ�= k��%�ෑ=���4��#o�;-;*�7����E���=�<���� zL���s�`���A.o�G�m�?��x�Mu�W���`moF˯�+)�H�f�M�&�����ϲ���6%�aj:�Mpp�}�(�-l̜	H��d˹�40<~�UxHj,��|��	��kޮ�Ԭ����}>p~z�r,,���9^-�I�~�џ0I� X�1��kޮ��g��� ��"aJ �!,|�8��5ǛHO��E��������~G����EX��dC$,\ͨ܉p����O,8�ݚ�Н�K�\7}�W,:S�.?<N��	�Ȓ�@{2귑�7��m�K�!�`�(i3+�uB;y�e����'�N��(���K�!�`�(i3I��
�[��b=��y��j��k����U{8�C,0�?��ʉ��%>�rG�<�]�Ե�����=�c�]�#+0�,��
������3bQ=�3�� �֤D�A��*ȑs;��|B���r����P�T��Y�"E&��� �
�V[Χ�>u�͙E��Q[AL��*���z˪�y��݈��0��JD����^C��}��3�zU�o�����L~΄gO�3�@�ɱ��w�.Y�[��թ�~X�|2;$�J�$�* a�N�ǁ�f�TpD��ZOUD�P�E6�k��q��־�W+��W�FwZNE�����A@�>�暩�͚+5�4��c�� D�_\���%>�rG6j�"Hs0vZ��ҹM�6(Mcg����*y}e!�|_@��0Ï�6]S*�N�ǁ�f�T��Ut>'L��nF���<�W�.�P�	��
�Q�}V;ƘdW��¹���e�J�Pn\���_*��I�Z�T�a��(ӈ���m�r����w�R���y�U��\JD>�o2��0v�6���P9d^\'@����y�w&�ŲVz��s�q@C�x�>���� �P��#��s�'	�?��[7�}�!��b!��u���j�4�<�..�4��un�H�@�#�rs�i��@�N3,(P�V��>'�o��&L*42�����`y���x��7��0��jOT���b�S]q�6��^�7s�9���o>��l%i�-@?d�s�8K,Q�\C䗬��O9�(UҔ����F����\/o['���Xw�j�7���ļަ��P݃��x���g��U-�e�P��|P��C>��ӚH�RtV�^��j�4�<�..�4��h��N�M�)n�w�'���b�'Beˌ�������)_�32����r����!�`�(i3!�`�(i3?Q�@X>#�t�{#	�x��>��',�$R�i�Yl-���{�G�!��A$�P������5d�Q'݀�=��`���φ��<�6��o�.�8�Hj\�����1:��\���F�`yx�>�+X�M?��y�!�`�(i3��@�z]���b��Bg��o���K7͍��|��W&":�ݚ�Н��T�T�y����O9�(UҔ����F��l_|�(K7͍��|��W&":�ݚ�Н�*qA����6\�4�@�� �-j�1tSjv�����l����� �'����u��r��!�`�(i3��j�4�<�..�4����%Թ+�O��b�S]O�lK�������[$R�i�Yl-1�*����"X��[A84Ы�"��m�q�/��]��V-[�ݚ�Н�;�x'_|~�RZ��P�k��!B>g����oo�}ߟ�r�Q�+���xҩ��ga@MxKkB)��5!�P�)��xuo��*lA�y�
M_r�>p�{C��Nq~o@G��-�HG($R�i�Yl-%�z(�~�:)�
�9��3�����ߤ�:C
#!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rG߸��S�Ȍ��7���9�:)�
�9�_����@�`���*1~��E�r�*��8lx��g�F�4�q�+ �Ǵw�T:~,�W�8"M��K���'���y��lD�k��k^�^)x�ݱ�5����`Ke4����F����,"��.J7h�4���>eC�r�&U������G|M�܊j��2�'���Xw�j�7��Z�qҪc����-W`9�,��R�cv�x�bIR�^Ƒ�Ӹ���p��j�4�<�..�4��� �I�8�Hj\��$�'�}�HL�U���WF*�L��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3K7͍��|��W&":�ݚ�Н�&�z���@h�D�-D���V5VM�d��a�c\���aR�!�`�(i3� 4� IkwqE1r-�erUڈ4�`,9�H�W��`�z��Y��),�B۸����H�V�7�}�!��w Xy�FZ?¤$O��P!3)T���t�f�2E��A_�u�N�ǁ�f�TpD��ZOU�_HĨ�ވ`���*1fĉ>99��;��|B������{\� C&���R�tG�"VA�ڦ�c4����,�ǰ'�J:��XD��/{j��W7�-ys᪐��*y}e�����2����Q�ʘ['Ӭ��yb5]��o�������Z��!�`�(i3�N��Q��ǺΕo�G�m�?���b�%ł�{_8�Y��=�}�Vݨ��}Dq�f�)�{6�U��w�.Y�[�GR�D^O@�s��M�t�3����mm���|��8�; ��8�Hj\��ň����L��b�S]O�lK��^?������X��O���r����!�`�(i3!�`�(i3,��G��z#�r��8ߞQ���l�N������d�Ѫ��O!�`�(i3
S�z�Q����h{��Y��),�B۸�ն�������N�����/ЁqVU��ס<�%�+���xҩ��ga@MxKkB)��5!�P�)��xuo��*lA�y�
M_g� ��9�C�;_�b�z'hۉ)��d�7�q�8��;Yv^����j�	l@ �&A�5C
2���Ks>�W�K7͍��|��W&":�ݚ�Н��k��M�vx=��X�&����������� ���J�C�M$���DФ���Z��!�`�(i3�r�+���ڳ������i7N�_H�A1m���C
2�񚡄�Ӹ�֧�5��,bXh��d���!i!�`�(i3w�.Y�[�GR�D^� #�~	�D�t�3������׻�!�`�(i3w�R���y�sL]~ц���X)Hp��Ɇ�5�HN��R��?�d���&�<�V�QK�}{�rD�W����#�!�`�(i3� 4� IkwqE1r-�erUڈ4�`,9�H�W��`�z��Y��),�B۸���Se���7�}�!��w Xy�FZ?¤$O��P!3)T���t�f�2E��A_�u�N�ǁ�f�TpD��ZOU�_HĨ�ވ`���*1fĉ>99��;��|B������{\� C&���R�tG�"VA�ڦ�c4����,�ǰ'�J:��XD��/{j�䰞��X"�y�.�g3Z�)V��B�1��b�vA#&��Q`���*1zY]�埅��!�ٞ�'�/��T;��%YM�	�v�3�x�y�Zgl�k�����Ղf>x�:	�W+��W�QS��:Z�7G��#{Ձ�=�niF=�xo�n���㬺����D�Ϩg��U-�e a⣃_B7�}�!����nސ�ѽv1a{J�����u_(�s<�L�K�������iA'R�	op|��G��}Dq�f�����,�ǰ��������2܌���!�QS��:Z�����n!�'��iF=�xo�R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#P��.J7h���/5U��nFW�JyS�N�*J�X�$����q(	�fI��)���W�w��fD�g�9��,Y��(c$�,I��)���W�w��fDbYގEV��2܌�)��/��;��|BMR��P.�IZƀ$�ֶ{�ӱ���9��;�R���5���T�}�@��'	�?��[�-���^�ߗ/�h.��t����~,�046dr����,�ǰ�X�t�q�6	�9ڈ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��
�V[Σ_[����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�����z�}�hP��Ÿ�v{7!I���6�{�Pe�E"��*X��[��7%^�W+��W�
�V[�t�H	�I1m��+o�Tku�����F�N~Y+��YR�7h�,b0V�u�Q�ݚ�Н���M��҃!3�X�뼥<7.���nH�W�f�?ǉ�=^�F��M֋)�[���6*bL�(Rp~z�r,,���9^-���2��̪U��֜��3�)ύ^��R�^Ƒ��f�?ǉ�=�����@���k�֩�4��#o��
�cc�V��ݚ�Н�W����vcy'��5��s,�ܠ'h|��W�Ty��5!�`�(i3�0�و�{s�ܱ?'�ފ�����x��7a�!�E�_�������� "5�]�/��@���Lt�2�t�&8�,������	�;�ݚ�Н�h�'f R!�`�(i3>N0Θ��ݚ�Н��ƿ�d���!�`�(i3M몴PBoT�ݚ�Н�?KYC'v�����S�Zq�%�V�m��s��d�?�+�p!�B�'��a� 7�J�[�_�C�6%���lи{K��i�g��C\�2x���?V��j�cZ)[���F�X;p`���v�<�$,�۞��	��P��J1zY]�埅؉��+�ْ��4F�;��%YM�	�v�3��C�M$���Xr��,��d���!i"(<K�'P��<�MP�`@���!����'d!�y]/�qF�ŝ��X��MM
��,=?�d���&��ݚ�Н�H���7Ә���|f����Q�یfw+�V��+O��cb>�g�D�fĉ>99��;��|B��D�$�eX����}�	76�&�;��|B���0�2uN;������]W&Z��E��3?�d���&�E=Խ����P�	�#�Y���I��� G�|]A��P�	�#�=��R-��#U#��F:җ�S��z���AZ���d���!i��9Ӌ�6Li��.��1�:�Ω�=A���>�LZ*IV��ӓ������~H	��`��,\ަ�It��+g[����=�-�o&l������g����=�tt"���O�����J��a�U"����N��Sx�M������p���,��2��������")d���ݚ�Н�Q١Ӿ�$������i��X;p`��ļަ��P'b�be`�t!�`�(i3ct�:��RE��]n��X&|a�#�I7��-5��5Z��=��]zŎd>&�&i�������kޮ��R�^Ƒ��f�?ǉ�=�B�6�N@���k��-��W����vcyj;��q,�zg��p����8��'@���k�� tZ�u���ߘ�)�Ij;��q,��z�_�Б����!�`�(i3�������a����"�$,\ͨ܉p����O,8�ݚ�Н�Gظ0�����@;w�$C,0�?��ʝ�hy��Q�#<4^�>N0Θ��ݚ�Н��ƿ�d�����&I���m�
��,!q�\E��0�����?Oǖqo�_����m6(\�]���f�?ǉ�=W����GS�*;q�j,���-�}s�Z�|�X[�m����!�`�(i3+�uB;y�L�6yd(�~��rͤ;��krk�ɍ���>Pҝ4��/��t]�<Lzg��<�=Lk��D5�|أͽgF"?�Q��ǺΕR'),��`�C,;�m�~�?�d���&�x��7��NmyM<�G�ۺ�Ub�!�V��u��i�_:�����k��$�8�B���ow_;O
�J��:����1�����j��G�m����t���[����<���/�sLXNAA�����}Dq�f�����,�ǰ����������^�)ߋ����-V��	��yG��Γf�-I�p��g�`ks�F���;_��8W�w��fDy�^ecK̅�8�:����	ڱr&�zbYގEV���{����/V��rU�w�⽒��8�>r&���nH�W��^�̷ؠJ��:����g������V���S����,vQQA�q�m�,�5�%]����8�B���ow_;O
�J��:����w�.Y�[�����V?�_.��45�$��cז�!�|_@��0,���1����,H/������,�ǰ���������{����/�_��.���9�Z�y�6nZ:ӄ��8�|����N!�֏^�M;�¬pX��D�P�E6�k��q��־�W+��W��r�+�����i�g��QZ���>�ĩk(�CQ��/5U���F�SRTpI��)���W�w��fD�g�9��,Y��(c$�,w�R���y���,!���f�|�H��4O��A�6!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc%�o�T�*9������ر0%W��2s�1��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcf����5�CX0��W@^H���%�#�o����q,� L���s��$�Z;��|Bq�D�7�P-7�vqq��R'cf���³5��*�7`����\Z��K��qb	��G��W+��W�ƻ�.=�+��T����oGo�Z�������/�)��ɖ`ۺ�����ݚ�Н�����S���� "5�]!�`�(i3A�sxW�O�Ji�];����R������y�����/��b��7<RnnB7Ԅ��W���`moF˯�+)�Ww��g�1�Z���=�,���9^-�L/���?T�x~1�@��@�Ce�<�˹�40<~�>b�eIG�5�}�]���p.0��I�![�Do�9�ݚ�Н�s 3�:��)�[���6�5�9�(��4V�����S�e����kn4@Q�/�!�`�(i3�G%�MP3��\�d1o�rs�i�CH����.n�Hb�2�Ǐ��Pn<���r��N�T ���t�=�v��*"3���'�C}ߦTd�n�g��U-�e��W�s���Hb�2�Ǐ��t��ۧ���Ɖ`���|�F����A�+�~@�\����F��aQ��T�\ ��B7Ԅ��١w��zj~�X����Z鎬�������(���VAD<��'�WdM4@�N��L+@���w�K�R he��as�C�G���-�p'�"�hPW���[f=HJ��n�eR���>��WdM4@�(%�(�Y+�(���B��U��0S���NB�D�u.?;�^H���"X��[O+oF��!�`�(i3r�x�e�X�	[F42���ON�C�ժ*)xJe�2��}���C�#�J�{H���7Әi��7u�`��Y��)����*�~p�R��M�!�`�(i33L�*}F��ߔWň���
�
��(:��IK��<3Lv	̅���X;p`�(�����
�:qEp �D�lh8t����s}�	76�&�;��|Bk�rOj��@T�J�E�w�R���y����C��CX0��W@^=��#̈́Ia2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!;:��t� �Y	��n1N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���X`
�2����1	�v{7!I���6�{�Pe�E"��*X��[��7%^�W+��W�}ϼ 8�����?�ؖt�_��<��d�٣���������ݹ�0�������P�I��RhF��K�X:��3j\	Ov��+���LQ���"X��[��Q[R�7���PM���KPkqy�{J�t��Mhm��+ r���7���?�_�#fr�L��ϸ��#|S������3[�u8�~6���q���)�� �t���������z��*�7`����\Z��K��l�`�
X�M�]V�H7'�R�^Ƒ��!�`�(i3��ߐ�*׿j�h�<��k�+9=8��ؤƼm��P���ݪ��	QY��K*�+W���F�^�Y�7#�xI���E���v:ι�Y+W���F�^�g�&�0m�X;p`����0/ܤ�(g��V(�G�&���k��,�:�N�*�x֭�h��Oo��0��7�X;p`�l.�	�C˟B�'��a��7��r�=�&8�,��Q�L��
�:qEp>c��?ӗ&8�,�g�Hn7�(��wӨj]h��_--���g�_�C�6%�m�;������/�sL�i��NU�q�\E��0</���/�u�k��rݾ(����C������Ce�*n�/a�~~��}H_��i�;��%YM,���4���I4��欱���j���u������>?�d���&�x��7�֎�ٕ��j�Txk^���%�>�?1�Z���=��#t:0���nS�3�ǻ��d���!i�q�9�ͭ��?�ؖtO��cb>�6|��ŌM�H���7Ә���|f��I�{�P�Յ.�g3ZrZ�0m�\���ٕ���E�i�m}66j�"Hs�l��J�&Dv��Y2\aT��3G?�d���&���H�ݵ���P�	�#���@F�_+�զ�����P�	�#�=��R-��#U#��F:җ�S��z���AZ���d���!i�%�_F�1�� ���J2��������������]9�(b���J��:����\o�LCd藀�)�_f����/�sL|�a;�{7s�9���on�-�6��
�jW��D���M���R'),��`ޔ5:�7�+p�i�_:�����k��$a(􆿳����^�����8-|�DSƏw0����n�k+}�I�?g�f �H�Z����dn��A�������M!�`�(i3�,\ަ�It��+g[�!�`�(i3��[<��	$e�7�3`�&8�,�뼥<7.��H�ʱˡFZd6�o�!�`�(i3w¹��<d���<
DN�!�`�(i3|�����ݪ���k�+9=�v:ι�Y+W���F�^�Y�7#�xIvє�&������0/�e��9�SW�Ty��5!�`�(i3�ܼ�Y�{ �=�%���]n���M��eh��y���b<$�O�媾k��M�k��,�:�N�*�x�/��@���Lt�2�t�&8�,������	�;�ݚ�Н�Y��
�iC!�`�(i3Tl�������l6������!�`�(i3�X;p`�YmC,igu�wӨj]h��_--���g�_�C�6%�m�;������/�sL|�a;�{f�?ǉ�=q�\E��0</���/�u�k��rݾ(����C�������|#HK���t]�<LzKj�`�|\{ف(�7���<��Y����}J�|���|���>�q;Rm�5�O�%E#P����&��t������~Ձ�=�nx��M���U����z~�ŝ��X��MM
��,=?�d���&��ݚ�Н��G�6\�堌S�����*��i7B��`	�K$$�������]���z2�T#��(�&���%>�rG6j�"Hs������r�r��HxjHN��R��?�d���&�zY]�埅�,Ǥ���(m�ڨ�hծ�.�g3Z�`�e�%R��	7?���x�;��XB$�6�Q��O�بeD�I�,����y���Z��Zt%��m&<��dn��A�9�2�L��f
t斃|�q�^"�HN��R��?�d���&�8>�"����ڻC�i�;��|B�}�+�㟝+0�,��
�䡷G�`]2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��o���sp%�LY�V�*�b֟�;���H΍䂌N g�}Ty�i <��m>OM�Ѫ r��F'�8c8Y=o�|`�,���;���N;������#Pר�xfa�X~��`�� ��t�ða�F��u��.t���xN�����@0�6�����S�@� �V�s�����%82���
qS��;�$M���g���w�*2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}��gj�ݬp+��T�����h�6ؖ[!�� Q鹈��fq�/5�����6��������֢&@��&����Kp&�@���k�֭AQ�0GȨ��_�\G��4�	B45j;��q,�i�ۑ ?�R��n��h
:h����c�u3���y��lD��,>��R��ӟ-����6%�a��Nm�ju�|`��P��a݃�j��C�`�/�t���E���� ������O�z���5$�<w����0)]��w�b^X�P��EގV�ڇ��t��˳3[�u8����ꀍ�@;w�$C,0�?����_F�k-�!�`�(i3���*[UxG���%>�rG�B�r�݇a�/!O�$-q�0c$�Zt%��m&<���_L�b�����Ee[u�;0�f�?ǉ�=r�x�e�X�k��rݾ(����C���h���?V��j�c�[N�&ѐǂ��%D�$o��)�ͳe��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�)� �~�K�����r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��"/���]�Q诤�e��C�`�/�t��cm�@�ᩖ%�!����5��fH�6J)�s���-�)��|���=f�}��U�����̾0���;���˔����vg�ĝ����a��X`��_/��;�y/Ә���@�ۻ|2���̂; ,@�� د<�l雲�fb�����m� D�@G��l��3\s��$�Z;��|Bc^���HP�a��t�'����9|s��^<4mB�@o��[�|�hJe�A>��*�X+��YR�7h�,b0V�u�Q�ݚ�Н��5���=\�B�wj$g8!�w� wk���,���9^-����y�,@���k���x�8�D"�����ׄ�R�
qtC�NI�Q4p�/Cj���C�1m�'*Gʯ7Պq�Y�.��x���"x�ś��5j�g��$P�M	�D�$ȨQ�?�Q,\ͨ܉p����O,8�ݚ�Н�h�'f R>N0Θ��ݚ�Н�Gظ0����t�%�Z?��<�ry^�%��C����\P�ʊQ�����J`�wӨj]h�vYv�������q��@����Mh?V��j�c�;J�*%n�+�uB;y��"Sek���6j�"Hs���%ˡ��V,b;�:��,����*���*-�,���O�]���N�����?�d���&�'3x)'�V�m7n,�
��W�.��A$�P������5d�������y�(����<m�r$ɓǃl[�Ƶ�1tSjv�?V��j�c3R�d�ܦdN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����}.z)yG��Hb� h�ҩ�?V��j�c3R�d�ܦ)�vL�����]W&fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vxI��S�ud��E�9K��;_��8W�w��fD|]η����Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9Y���&���'܍|Cy���QJ�wk����\����|ݔ�3�(n�'�(�S��)��R�^Ƒ��;��|BEΟ��
�U�a�(��^GѬ�_���t�T��?E-h��`f���sC>��ӚH�RtV�^�'ž1�|�'����u��r��q�\E��04>^!b!4b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3��Nh�=f[���������<�.�����8��GM��-����!�`�(i3�v�Wס���G�K$x/��&���PC-��i0Q�͹�Ɩ,�b�R؅�!�`�(i3q�\E��0����G�t���m�� �ݪ���CyW�f�tR�wX��!�`�(i3��Ě�����}Dq�f��3��C���H�� �YߥթD�[*�Bi�v�V���;AD�e�{�W!�`�(i32+5�"�����-P��F����~�;2V-W��	c@�^ k�R�e�0���m�e#e>�=�^݊<���He�ylB��-t���m�� �ݪ�򈟕��+�v�7��]�ݚ�Н�3��0����g����F����~�;2V-W��	c@�^ k�R�e�0���m�e#e>�=�^݊����xQ�e�ylB��-t���m�� �ݪ�򈟕��+�v��t���?�� h�ҩ�!�`�(i3�lTN��I���q�}���{BO���5�%]���a(􆿳����^��!�`�(i3��jVѭ@!�`�(i3u?�:�H�jsrCm�k�J��6�d�t��w��X�'����u��r��!�`�(i3q�\E��0��@Z���rs�i�}�O��LTSG��ʎ�=U9��R�^Ƒ�Ӆ��I�ѪtR�^Ƒ�ӆ�v�9��!�`�(i3�����!�`�(i3�wӨj]h�(%����Z鎬�������(���/%Z�ڄ^1��#ƌ/B�ݪ��2�r5�����jV�{+�fbmDF�!�`�(i3���%>�rGO�D mWN!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ o�n�J-�ƪe�0c�)�Ul����,�ǰ	r�R��Z����i�|7��_	�s�t�{���6������]'m���G�K$xE�p4rqG7]u��
�3�R�^Ƒ��;��|BEΟ��
�U�a�(��$��,Ix�6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3e�v��ҵl�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r��pT/�GS��%�����d��-��![L��^C�+a��o���H�RtV�^q�\E��0��@Z���rs�i�@24b��H�[���wkL�1p/-��G�<6�U����z~)���	6�
�:qEp�;�P�t�5fĉ>99��A0ok�׹�3��܌o��oŵE=��X�z��V��	��y�߬9�6ש`/V`L�v*2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc� ���j���Gɾ>�z����5Y��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�Y�Eat2�\��n�q�����"?��A$�P������5d��n4s1��7�癆cgQw�c4~Nr_�mS8<�n��!�3�
䖬n���/ ���we��0�U+�qbp@���{$@d9mh��n�tr�yÊ��_
�u}%GP����ZLN�	��� [-�9����G�^��D��!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^�wg�]��l�
@\�nQ�rV��q�t7��-����!�`�(i3�d�@���GU�lP4��/����*Q!�`�(i31���~�>=���#䖬n��؂�nF���<�W�.�P�	��
�Q�}HN��R��bP�63Z�t�G:w���he���!�T�1tSjv��>=���#��he�վɢ���he�U10���i!�`�(i31���~�>=���#��he�վɢ�F}���V6M��C��]��ġ��,���t+X�}��NۥUn��g��� �:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�J	���/a���Q=	+�{�*��{�ՖR���D�8�����t�T��?E-h��`f���sd=��¾ȼ\���F�`yx�>�+X�M?��yЃt����}����˃�I/ ���we��0�U+�qbp@��t����}�H_��#�Ր��V��e��0�U+�qbp@��t����}�H_��#�������i�e��0�U+�qbp@��t����}�H_��#�՚`��n����{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^Us��K���(yJ+��ʤ����3�W���b�0�T9��JG��NۥUn�+
�Tn@H�oi���:�l�^���;�jmT�#�>k�N��^��hJL��;���N0�!5R�u��r��;�jmT�#�����3�Ⱥ;
J��0�=<MW�-}�	mp5���%�+� h�ҩΪ���l���oi���:��*�·Op�r~�h��ݚ�Н���w�w:�!�`�(i3T9��JG��Bf����{_8�Y��=�}�Vݨ��}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t�Zj���
�d�@���G����B� �b��!�`�(i3�D���s����NۥUn��5��\���� h�ҩΪ���l���oi���:?�Bo���],��%s��'��_sN�">�������Ra])n#���r�����t����}�H_��#���վɢ�F}���V6��%��@qf���-A�¤�x.�Knqrh#��Y�
9mh��n$��k��3��,H/�����%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��jϤ�Lǀ�r4��3m��Jw��3�+=�4o���+��+}�K=���e���Օ��qvdЧ^{�jM|�"D5�O�%E#P��=m緒1d�;q3�)�U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩΟ/��mS%y�W�CbE�{_8�Y��=�}�Vݨ��}Dq�f�	�)��&ghRV��RK7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv��B�'��a�S���%��������f��1.X!�`�(i3;d��'�XƤ5_���H(�T�O��{Tɀ�"'��&އ�[t�Y81�d�@���G�X���.��ġ��,H�Ћ�r�H�RtV�^;�jmT�#�YN
��)e���^b�~H����8�O�5���1tSjv�!�`�(i3�/��mS%�r\���%����g\>������
�:qEp'{w#/ B!�`�(i3	�)��&gha�E�Rq���my$�N��o�/���;!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vxK���q
�&�lV*�]�aT��3G?�d���&���#��� �Rɫ�%�'�M��+��+}�K=���e���Օ��qvdЧ^{�jmWᅫw�5�O�%E#P	�)��&gh���(A�,"�(-w��N|;��|Bʦ?�H#F`�� �R�!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcۖh��)������E��㕷�f�Ux�_����+�b��T�Q5�r#�.�O 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �3 �����|��sQ�G�=�_�7V�o��_�Rv�䩲$��8��I�:Fa�7���z��O�|��/7*f'�|��bs��2[�a��o���H�RtV�^ϟ��7�4ÿ����Ԃ�nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r���Zj���
],��%s��ԏ ���ԭ�m��3��p���H���6Sa쎑t2�������50f
V��.ᬵy���Ÿ�`u�1tSjv�V�Ո��+5�4��c{�"�S��+�ϸ�i���U������՝� s�#���k$ ,��G��zł)w����ۥ�Y�mK7͍��|��W&":�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�������ł)w�����Al+�HB�����������mA�ѕf�f�_T:5�����2������}W`�J$˄���Z�׭ �k�3���u`�`�A ���\��o��_�Rv�䩲$��GQЌJ
��`���φ��<�6��ڱI�̘'np>�#�=�|#HK��A(�c���_G��Hb� h�ҩ�9�{�Jj3Ř�z��l �vPu06��K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv�V�Ո��+5�4��c��W����W�/�#+*f|��sQ�G���+����rV���qޤos�em��ܑ��y���8���/�DY�7f�P:��z��l J	ibP�v
�:qEp�;�P�t�5fĉ>99��A0ok�׹���C���N�ky�A�掲t m^1r����,�ǰV6f����np>�#�=���-Q�OP���N��-��f���]_q�g�]@n_���?3Cy����]E;��|B����UrV���qޤ%�n#� �nF����bS��jarV���qޤܡ��F؝=��/z*x�n;��|Bs�'��OWnp>�#�=��Al+�H������B��/�����x��+�]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7N2��j������mA�7�癆cgQw�c4~Nr_�mS8<�n���*y}ep8@)y@dl�SB%��I97��EN�h�h�u+��.ᬵy���ܝi���ؼ
���$����G��s��c�,��G��zB��/�����I(����K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н�`)[�-hnhG�W�W�/�#+*fG9�:Q����t[�L�a\Y����+���LQ���"X��[��Q[R�7;�jmT�#~��F�����������yN��7��aq����i��oZ O\������U�._�nQ�rV��q�t7�l��8����aGl��Z����pG�p�P>M_���u��r��;�jmT�#`)[�-hn���+}ȵ�v��ONH!�`�(i3����ҧG9�:Q��� ɦ���AԢ�a\�Zx�.����#��o�TX5Ȭ7�j�W����^��D�Ϝ�}Dq�f��	��x��ݚ�Н�,��G��zB��/������R�s=Tu��H���9�-�a��W|!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�ȌM��:�3��H���9�4���qB�Kj2�K����S�p�$@PJ+5����E�EG9�:Q���OLF+Q�>	#4�a��?b�@</�P����B��/�����>���Si9�i���>6�b NK�+���w� �~�^h�	�i^䖬n���n��y��a3}PR�]C$�.9�?	���58���d�@���G^?������X��O���r����!�`�(i3!�`�(i3����}>Y�&�-���k%�B��;���N���%�K�W/S��8(�E���Kt�emW��EG��-WBgW�6�h�g+�{�*,���H�z��ݠ�s����J��ͻ����8��Օ��qvdЧ^{�jmWᅫw�5�O�%E#P/Q]=��7�k]m��&k@C�Ɨ0z�cULj� 1�B��/����9-��g���t�
�:�WdM4@�r)1;�Os�rs�i��5O
T���ihc�ؓ;)Ve��˅�D�����R�`�|��K�z���k��$a(􆿳�3�m�
2]�����,�ǰ	M,��rER��p12���v1a{J�Զ �3 �����}c��ko#1^���E��'Z*)�?�R��nj��P_Q����t�h��W+��W�����"�>�3�eZ~��!���c�A�L'��B9[��EF�*���]�!��	Ǹ�y85���Ü�ۯm&����T��V��l/�#>6�b N>�3�eZ~��!���c�A�L'��B9[�o6Z^p�'���Xw�j�7��>6�b NK�+���w�(�)��c1�a-���7a
��r��L;Л����:<��j�.�g3Zv���� �_a���zz�2[QvA��q�q�ʩ)!��w������"��d���m��+�Z����y�+��Y����S���� "5�]¥������]n��-��A$�ʁ�bDT8!�9 ��h��ˎ�){�Ysy�t��P$u��&8�,�oa�}��p�-�o%�'b�be`�t�D�&��� �4V�H�%p"��RR,���D�#��-�Vgh�䊉��	��J�6p�N��2��,Wc��I�W�"�Ů7�6��,�ݜt��ϑ_�������� "5�]3Lv	̅���X;p`�(�������0�&�ͭ�U젩`#�4>?� �1%��C����\P�ʊQ:��IK��<��_(x��`�:��]]t}c��ko#@�jw\�D�wP�/�w�I7�w���c�ۡ��T�
jl��.�t�r�$6��y�H��}VV��5l+��@-�-'͏��������FG�n��,\ަ�It��+g[���x��&^�B�wj$g�X;p`�>6�b N�A�7�dA��L1�l$Q
ˋ!E\1�1�ҕ-����s�;�9�����:�.�Z�%P{����8��T�h���}둮j\����C$L$E�͆عE���ؼ($��:�e�hfH'��!�i����VZDf�?ǉ�=�2*Q=F���q/���<�����7
��+qѭ�+g[��_F�k-��苇��Fe#OOJd֯̇i�d�?�4�0 L?�p���@Z��9��稕�a�/!O�f�?ǉ�=扈�N̮�$�WdM4@������p�n���:��]]t[��m�UAIYT� �?��	`��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcۖh��)������E��㕷�f�Ux���蹒��yb��T�Q5�r#�.�O 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��Ɔ ���ڣ��>7�v�\�b͐�	}�@�r�<Uee���R�}vJ^j���W���?�d���&�db�\EX�b�'Be������>���$���gE�s@��b�'BeXxg�H�������,�ǰ���9kn��회�h�#5���u(_r�r+���U��3��aO�R�[5C�R'cf���L���BN�.ᬵy���9��Pሐ���Z���G�dE�h�k]m���1��̍눸�)I97��EN��()��#u� �GR��shbvk~�#xǩ"�4s2Zx�.����#��0�8�ڇ5�[�x�X���+���LQ�g}|�H�/�����sc�̆�!Yx�����!��,�j:&AԢ�a\�!;���}�ߜ�*�l8�b(�����-\71v�<om��-T�"�N�i;��#��F�r�f�tm�;�������,�ǰ���9kn��회�h�#5�5�s�p p2���i��_A���e�6|����_	��[���R���P��J-��;qjl���j�ވz:u�,䅽�~TX��MUǪ�^Z�e��1q��U��)���Y;e�iK!���d.���+�^n=\f�5>��YL�P��tõ���lF���d H���� �'ž1�|�'����u��r��W����G�iA'R�	)m��p���+Az�q��{_8�Y��=�}�Vݨ��}Dq�f��Ɔ �����O�����C�1�r5��(ә��nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r���G�dE�h�k]m��F���d H��(ә������D�v1a{J�l����Ȃ���C.�uW���ٸ��N=�z��S)��.J7h��C�x!�H���J��Ӊ�,�O�%p�+Az�q�N��	�Ȓ{A�dha#4\�0l�sf�e�}s�P�g�7�M^���H�L���%>�rGO�D mWN��Ě���aT��3G�IX0F�M��&Y��V�f�\�`"(N����ʴ5�S�H͞ {��b�'Bef�Ϡ���N��	�Ȓ{A�dha#4����ʴ5�����d)�z�~I�x�H_��#����Y��<�;-;*�7�����G3҇
N��	�Ȓ�cЉ�M�@�\��?��b�'Beͧ��&�~LI���p�����d)�z�~I�x�H_��#��jnbAo�[�x�X���+���LQ�<��N�ܷQ�,!���vc|�M��8�1�:�Ω�����|"#fr�L�t�iZ]XF�hx��G��N����p$��<
DN͗&8�,�nU�gF�r�f�t���MK�L��.��֞�������i�4��%�;��g��cH�wA�?�D�g��ۤ���ֻ���~��a[/������N�� �ȳT�_�O�0Pa!�����V�`�4G&��z�D�&��� �4V�H�%p"��RR,���D�#��-�Vgh�䊉��	��J�6p�N��2��,Wc��I�W�"�Ů7�6��,�ݜt��ϑ_�������� "5�]3Lv	̅���X;p`�(�������0�&�ͭ�U젩`#�4>?� �1%��C����\P�ʊQ:��IK��<��_(x��`g�%Y��̗0z�cUL#������b�'BeWh4:z�]MD�wP�/�wK��=�C�b�'BeXxg�H���M? D����j��=��
�lo3��$����'HY-��
�C�Ʌ��HW�ǳN8�e���x�l��1�V�ܡ���¥������]n��-��݁.�q�0��E|�,���E򾚲-/E8�)�[���6�X;p`�g�]@n_���?3�B�=9ODۤ���ֻ���~��a[/������N�� �ȳT�_�O�0Pa!�����V�`�4G&��z���Fz�^P��:w0I� X�1�;LV^Š�r��Lo�_���Fz��2*Q=F�k�mD#V�C���b7O�4�xKKوx����y���ݫ�ф'����2�_�������R#���:B�V`ЪF�,�U6>���|Z�,:g�.X:$����z�����	�;ׇӭ����"����M몴PBoTׇӭ�ш�_(x��`g�%Y��̗0z�cUL#������b�'BeC���YXA���Fz�@ E����]�;���Vнv1a{J�F֢O܋^����R��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�-I	�\�'��i���~�߅��n������������ر0%W��,��l�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �˥�'ܤ",1u�#+�����đ��%�/��Z>LUc�f+�Vr���F�!��c�)���A7��!=BM��~X��ͷ(�-[BݭsF��Pg�ÿ������U��)���Y;e�iK!���d.���+�^n=\f�5>���ah��ol�~{�Žxjzӝ���I(͂��-��������ҧ|���|��i1.��2�8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&rG��Hb� h�ҩοa��=����
�
��(-�y��j��T�B�X
��j��8�u�ׇӭ�ѿa��=����
�
��(�h �g��M�&�^���RD§B ����z�le5W�F�h��
�
��(�h �g��M�&�^���ݵ�Q�n��T�\ ��v��؄aX�,��G��z�T�B�X
�*��U�-��>&'�5�M�&�^�������W�HN��R��bP�63Z�t�5ߧE4��Fr��j�@�f�smy�Fu^��0�M�&�^�������4��;��Z{oBQ��;��O�"������$���(��g.Cf���ϟ
B� �r�_�B&��p��ѿ)�L&�Fڱ���E�-�o%�烒�]������B��/Nߜ�*�l8�b(������l__��S1�c���Q��ǺΕR��ӟ-��G����JVW{�-v���m��3��p���H������7Pr��ġ��,;�4q"�?�d���&���>�9�=U�d�#�b_�MN�8C��D9�C3x�В&=�y�q}��:��)gi����S���� "5�]�D:���@���k��!�`�(i3��4��#o�;-;*�7����E����){�Ysy�t��P$u��&8�,����揺hvl��9�h �=������-�S�h �=�*�a"4̥�0�L�p~z�r,��:fۇ�0�=<MW�-}�	mp,��_А#�<om���Ϻ� ��H����8�(����������cɧ �GR��shbvk~�#x ��M��.ᬵy���-�ki�;Q�ݚ�Н�ss2����
)\Y�����'u���ɿJ��ݚ�Н��W�"�Ů7��B����3�=���!�`�(i3�2*Q=F���q/���<�����7
�e����kn4@Q�/�!�`�(i3k/�z�xEQ���*[UxG!�`�(i3���ꀍ�˺�Q���f�?ǉ�=��9��稕�a�/!O�f�?ǉ�= �@��&}��s�H��rs�i��='̹Z�;�C�x!�H�����j??V��j�c�;J�*%n�fePh����$q6�E�5j��/z*q+6j�"HsF�prB/ˬ8��� ��K���.v��>oKk�����jֈ�U�d�#�b�.�lo��y>'MM귈nIg�R�5��/dV�ļަ��P���]6����(����c�n�R�HM���#g�8����f���-A�¤�x.�Knq���;W��ZLN�	���M�X�FG�p�P�➁q��H�g 6ͥk�0�=<MW�-}�	mp,��_А#�<om��������oK?�d���&���>�9�=U�d�#�b��Z���Y�{'%s��jb�ܳ�/�����up�͸yob����,�ǰ����x0�J2�*���fePh����{׌ISU�d����\�a���GE���T��>����$R��׮	��48ܼ�P��������.�5U2��53��N����"�|j~�]�������:�.�{4\�������Fp7�D�_�k�W�A�&hH\�LZ:�\�Ԋ�{Tɀ�$����nQ�rV~��s�N�h�5,Wlr�r%)cAS�|Gv������9�f���-A�¤�x.�Knq���;W��ZLN�	��<ϩez
����Z�ׂcO%��PR�k`���)��b%B�@o��[^�}� u��=��5W_~H	��`��,\ަ�It��+g[�N����p$��<
DN͗&8�,�nU�gF�r�f�t���MK�L$Q
ˋ!E\1�1�ҕ-��vؾ���D�_�k�W�A�&hH\#j~X�6W�A�&hH\���2*CA>0�1ۍ�h �=�Y�Eb�3��;�WQ�.p�2������}u��Kh���m��3��p���H������7Pr��ġ��,ˌ�����'�̗����Qnջ�%�f4�����p���yN��7��aq��G�n���t�;���N�竿��c�/-�Q�����4��)+�[Z����&�+x��z�@CP&Aq2Y��kک�x����y�mZH֫&��5�q	�jo�����<o���D�噸��\i�s�h?���+qѭ�+g[���hy�NzK�}TR��b=��y��j��k
e�3+{�i�m�T��!�`�(i3&��s���qz�Gb��P�!�`�(i3扈�0��"��S8�vV�y��F�k]m���~�þ�w�wӨj]h����dЕi�����,t����3dТ���S֜���,�ǰ�98#.�Ƌ�Z{oBQ���|�D��Yi���t�E��j�AkUx���6`������Ԁ"<�h^�hvl��9�h �=������-�S�h �=�*�a"4̥�0�L�p~z�r,�d�a�{u�䫟۟�>'�o��&L��)��")�0�=<MW�-}�	mp,��_А#�<om���Ϻ� ��H����8�(����������cɧ �GR��shbvk~�#x ��M��.ᬵy�����	��u a⣃_B�h���Q�kUx���6A
�ߠHZ鎬�������(���'�jh�,�cЉ�M��E�
��6j�"Hs�!Z#bl)IA����Cj����tLWa��U�@����ц�2CW����+�]E�]��q�}�ٳG���|U���X�[⺁�zfePh�������	~rV8C��D9�C3x�В&=�y�q}��&��z lc�x�l��1:�N�*�x:��+���������i��@�����[�x�X���+���LQ�f�?ǉ�=�gCu(o?C!�`�(i3uwТ�
2������}-c5����;�WQ�.p�2������}��T�� v�0�=<MW�-}�	mp@�s�p���.ᬵy��H0@&ɡ��Օ��qvdЧ^{�ja����ȓM�Me��U�3B�L���_��VP��{˒��Ύo^ZK)
�����-VL�k��V��6:�H�?Pc�L�x·I3o���<�6�Q=L�УΛ
V�x�:�	͛���b���4��)+�[Z����&�+x��z�@CP&Aq�K�^��Q��G�S>\.�!::tm�0�i.�9�O�G?X2�K��2WI'�=��y0��s���4@Q�/���hy�NzK�}TR��b=���|��p��PIQ#�C,0�?����6[��u�9k�\,���m�
��,! �@��&}��s�H��rs�i��='̹Z�;�C�x!�H�����j?{k�h�+�>��y��j����tL�YK4U)	�����ц�2CW����+�]E�]��q�}�ٳG���|U���X�[⺁�zfePh�����|υ�Ffw딶�<?�3x�В&=�y�q}��&��z lc�x�l��1:�N�*�x:��+���������i��@�����[�x�X���+���LQ�f�?ǉ�=�gCu(o?C!�`�(i3�m2��W�����}>p~z�r,E(7j�������}>p~z�r,���)�b�2������}w⵾k���yN��7��aq��hx��t�#���F�`�ã��Օ��qvdЧ^{�jb&P�"NE�<�6�Q=�	���c���KT
;��b�^"Bɨ �����V��m5Y)14 (�C0��٢�[.\�G]}�$C��� л�t�|̸9�73A}p��)�D�&��� �4V�H�%p"��RR,���D�#��-�Vgh�䊉��	��J�6p�N��2��,Wc��I�W�"�Ů7�6��,�ݜt��ϑ_�������� "5�]3Lv	̅���X;p`�(�������0�&�ͭ�U젩`#�4>?� �1%��C����\P�ʊQ:��IK��<��_(x��`g�%Y��̗0z�cUL#������b�'BeC���YXA�2��}���zgm##����Н���A�Y��|Dvܔ!�p�F�`n��i������+Z}͐�	}�@�r�<Uee�N�����$��̼�K���Z�׭ �k�3I$T�w�����+!�/}�u�F8O*�E`��f�A���yN��7��aq��hx��t�#���FӪ�c�g<;��|B�V���pu����p�5�"��[�B xh`�@�7�^E4+у��b�Bϱ�]h�(NAP/i�\	t�R��-�g� �GR��shbvk~�#x�l7�l�r�#���F��|}�&��3���.1t΀�+I@Lv�@[�JJ1��P�M��j�)6)-
3���WS=+E�
*��H+2siŞ�W�%3AԢ�a\�h�_e�8�4sg��ǎ�*��Zۉ�L�溥����v�8:hJ�tV�nQ�rV~��s�N�$²�ؗ$_Krt��qc�~�`롎q�C�r�X8g��mT�Of���-A�¤�x.�Knq��H�����ġ��,a��bt�eC�����m�������y	����F��،!|�α+s���s�֩h6$A����U��)���Y;e�iK!���d.[�����(����<m���"sS<�0�zG�������&G!�`�(i3v���,Ͽ�2[QvA�ͧ��&�~L~l�d����!���c�A�L'W»��`�{B�P��w(�f�� l��}I�?d�G5V������yN��7��aq��͹��e�[�.ᬵy����{!�)X+J��a�_݄:�fnp7Syv�Jы�^�)w������e��)��{}��M�+�'�̗������*��fPP!�`�(i3RnQ���_A}c��ko#)Ӄ�X��~l�d����!���c�A�L'W»��`�{B�P��w(�f�� l��}I�?d�G5V������yN��7��aq��͹��e�[�.ᬵy����{!�)X+J��a����P�L�E��w*��@�1�˓:�B��>Pi(���B���Q��ǺΕR��ӟ-����q���Ĺ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3܌;���d��-��!i��$>�cQ׆��p0�Ĝ(�IyI�1"��f�Q׆��p0�Ĝ(�IyI�(�����'����u��r��!�`�(i3J���ٯHb�v��ONH!�`�(i3m�����Gd��}U؄�k]m�����m;
h�����B]�Pd��}U؄�k]m�����m;
h���^/�M2!�`�(i3z��-��g���k$ ���y��lDR�6؄���c�ۡ��F</h,��.�W	̷_��yC��S8����2Ho��@��@R�^8�*w��T��v�9��!�`�(i3
������}Dq�f�;�jmT�#P"G�wk��g�e��C�b�g����P�|T
�ʪܟ��[�x�X���+���LQ��B� �b��!�`�(i3�H����AԢ�a\�ۯ���@Z�2[QvA�ͧ��&�~L��X��� ��Cѻ�~���e�)qP@L0��U���(�犽{Tɀ�$����J�	�LÆ��S1�c������b5�2<B�!yf�� l����jA��L�L�溥����v�8:hJ�tV�nQ�rV~��s�N�$²�ؗ$_�#,���R�u��r��!�`�(i3��k�C�-�<�ao����O����8Q������51�X�c�rs�i� S�xSVe8��/��u@hy�`�w��v1a{J��\>Pq������^�L��,H/��!�`�(i3�����!�`�(i3�q�9�ͭhy�`�w��v1a{J��\>Pq�������B]�PZ鎬�������(���Y�&�-�yr�/ӶWȶ���/�Z�k�ʆ-�(i�pY%���m��3��p���H����HRCJ��<om���o�p��F��0,5 .�U%{.�V#?p�&���A �80D� �Y�]��`�E(���B���Q��ǺΕR��ӟ-����q����!�`�(i3��Ě�����}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rG߸��S�Ȍ�M5b�&:|����*دHN��R��?�d���&�/�M�í��{_xGSn�����z����b�p����ī�����bL�'���IX0F�MV�ҁGG`5:�����+�^n=\f�5>�������Vmm�TF-���?4���R;�|#HK��A(�c���_G��Hb� h�ҩ�%��C���Q׆��p0~�5�H5m�v�&�k���������|e"%��C���Q׆��p0~�5�H������I*�&�v��/��kOT��ɕ�eYl�x���
��e���F7�Gh���l��,+)P<�ܓ�Y��+�t2�����dz����NR�p��@���|2Z��|��� �ҋ�;��}Dq�f��L�����B��2�k1�h�H��*��;�Â���ESҩ/��kOT١w��zj�X�X�>M�a���;}`O�k�4�����ˈ��`�@�./��kOT١w��zj�X�X�񳱅���^����z�嫋�T����|e"*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3&aD�4�X�X�[RP� .��ɒ�F��kB�t�x���@~H��k]m�����G�5����@~H��k]m���@� �
,9*�����
�:qEpNh���W<˥�'ܤ",�X�G[���7���B�t�x���@~H��k]m��E7�y�PjNh���W<˥�'ܤ",��E� ����e���,o�ݚ�Н�%��C���Q׆��p0~�5�HRoP��e�*�&�v��v�A�
^^3�V�C��k�HvL)��E��PT�Q׆��p0�Ĝ(�IyI�1������w5���iѹ�+�t2�����dz����NR�p��@���|2Z��|�����:l��0�5G,��Gc#����a4����dz����NR�p������jp����a�)�1�׀�<�6�Q==z!
���-�F�i��|�Uk�rDp!!v*!���K�5OoL!���}/
;$�Z��"�Y�<�SЮ!�`�(i3�L�����B��2�k1�h�H��*��;�Â���ESҩq���3��`��R�`K��"���վc7t��B��2�k1�h�H��*L]�f��e��
&YY��!�`�(i3g�>x�����H��6��b�4ƭ,�t��2� �צ�L��^�뢗�˯��Wނo̒.�9�lA�J�����١w��zj�X�X�>M�a���;}`O�k�4�����ˈ��`�@�.R��ak����`T�ҩ�	r�s�"���A���3A�n�+�sQ}b`�����E���v�RK��h�~s�K���Q\� C&����q��Z���Y�eF@�Af8�ٕ��(�W%����`ɊP�oT�L�ݚ�Н�?�C�KQ]˥�'ܤ",��Gc#�����O8��vW���V�C��k��38�h�3&���JT��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;��Ɨy�"c�z�
7!dB�c���Dx<�f�8ݵn����`Q�����^��h6$A����U��)���Y;e�iK!���d.O.C�U��B��-� �ѕC?"p���h����1�sH�RtV�^�'ž1�|�'����u��r��N
������Y�U��3Y��P4 �<�5Ɂ7dN�<@Iv��nt=:��:5A��pG� �l
s�M��KJ#�	g�˿��ji����{_8�Y��=�}�Vݨ��}Dq�f��L���������h\�L�O�c���ESҩK7͍��|��W&":�ݚ�Н��V��G F��x�⢄1@aw5�=Â��'e��0�U+�qbp@�!�`�(i3o� c �R�%1���%��K��>Pn��>�my$�N��o�/���;�B�'��a�'�7��E*��0U8��v��*����x����E2b�z'hۉ)��d�7�qĘV�52SG�U��@atA�ᴽ����rv:��q9+t�}�ݚ�Н��V��G !]�~F��A�mi�K�7�����//�ƍ2���lę�k�C�-�<�ao��6���z�S�yC�wbN�dN�<@Iv��nt=:��:5A��p�e�<Q��Y#ѥhZiC�������;q�{_8�Y��=�}�Vݨ��}Dq�f�I&!y'}�}c��ko#ƌ0Q_,�I����~uK7͍��|��W&":�ݚ�Н�^)�G�B�+�WdM4@����[y�K�/ ���we��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���d��-��!i��$>�cQ׆��p0~�5�H������I�I�߷�c/��-����!�`�(i3����6`X�/m>8Φ�ʽP�Rܷઍ����:~�Y����.��������h�4��=y����͘6��q��kUx���63��<�����ݚ�Н�G� �l
s�M��KJ#�	g�˿��ji����V��G �pȌ���]���E:�qL��n��p��b�Bϱ�fePh�����yf sg���}Dq�f�L��/\��=2���H��̣��O�˰�]q8k��.ͥ�H�RtV�^��.J7h����ly�P�r��n�Ŀh$�*�]�`�,\��ݝۺ���r��������]�Y�_�H��!�`�(i3�����!�`�(i3/w1z��ӊx�D�Re|����xت�����:~�Y���Wql����BM"���}Dq�f�HN��R��bP�63Z�t�V�52SG�U��@atA�ᴽ����rv:��
w�	������9�~�gz��8�,�@�VҒm�L��@�a��Hb�2�Ǐ��Pn<���@���(9[���G�������+��<�ao���#!��H�ȯղ!�`�(i3v���,Ͽ�2[QvA����[y�K�Q����!��Hb�2�Ǐ��Pn<��!�w(�y?fĉ>99��A0ok���H�����Yu���*Y��b"Wfי�b����{�6�o� c ��f� .):_�mS8<�n�ݚ�Н�t�R!ME��ߦ?�~F��C~/*�t�2�q㬑u����p�5�"��[�B���p�8����Q����.��$���g�e��t����3��v�9�ʘV�52SG�U��@at3Y��P4v��*�����*�R���Amr��8On9�*�����C.�u�X��I�ՠ�w�O�����|�D���H���~�����l���X�� QT��0+��?�DEu�>��-��4�1tSjv�!�`�(i3af��pD�Ї�6~��Ȕж�{�7�^E4+у��b�Bϱ�����ס�07Syv�Jы�^�)�:5A��p�Ra])n#���r������.J7h����ly�P�r��n�Ŀht�2�q㬑u����p��8��V\⯜�'�,LF!�w(�y?
�:qEp�;�P�t�5!�`�(i3�V��G !]�~F��A�mi�K�7�_�R��U��@atA�ᴽ�R܀{�!�`�(i3^)�G�B�+�WdM4@�%ρ��r�}6�/S� 8��/��u@�n�Jt�g�v1a{J����w �!�`�(i3I&!y'}�[��m�Uƌ0Q_,DE(_
/�n�Jt�g�v1a{J��A&��R�����%>�rGE�}�Wk�m�ڨ�hծHN��R��bP�63Z�t��ܐ�}Ď���!�+����=@�Hhg� آP��n~���=2���H��̣�� �<�5Ɂ7^���H> ���8ѳʳAM��KJ#�	g��7������Hb�2�Ǐ��Pn<����5��-�����dz����NR�p��@���|2Z��|���-��4�%m�Y$� 1Q#�6q�U��@atA�ᴽ�t�2�q㬑�M�{�|L��!ߩ��`4%�fZF�Gck��x������=l�H���3���� �����G��D�h��y@�Af8�ٕ��(�W�5���^�.I�����wl53�e�%^oe�Y���q��w�X�X�񳱅��5��]���h��N�M��z3:��K�z{�� ��C~/*��f� .):����6`X�/m>8Φ�ck��x�����ٷu�/��kOT�n���h�n�&Sq�a;Uйc�e�0�RAL�!hy�`�w��v1a{J��]%���0��8ѳʳA���9�~��� �������xNetҌ5`��K7͍��|��W&":��u[���ew���m����x��O rQ��qD���FD>�v��Pn<���S�׫�hc�!ߩ��`��0+��?l�/��X��MV�,oF*�L��!�`�(i3!�`�(i3!�`�(i3�q�]��~S��b�Bϱ��Y�X-�jjL�E��w*�8.����6_f.�}�ٷ/Tu����W`GU�!i&G�\��u���9�9��g"c{r�Va�irR��ak����`T1�h�H��*�������fF*�L��!�`�(i3!�`�(i3!�`�(i3k��_� ��(ӈ���l4Z�/��m�$����F�f�J��K��>P�a��]�/֢��s�Kȓ�FG���<���+tx�D�Re|����xؑ@�VҒm͏ڹ�)�u="��x8I�t�2�q㬑��&g�hh\�F�u������ހ�af��pD�Ї�6~��Ȕж�{�7���LM��Q�&�-�8Q�F���"�>mS@*�1�:�Ω�����|"#fr�L��ϸ��#|S������3[�u8�����$G⃍�������Z�N�j��>E�%��*d��:=�;�.x9�S{�$Q
ˋ!E\1�1�ҕ-����H(�T�O��{Tɀ���S�<Ԣ�E,�J�|R�ZLN�	�������^����8��T�h���}둮j\����C$L$E�͆عE���ؼ(�K�^��Q��G�S>\.�!::tm�0�i.�9gh�䊉�䞘gx�n�W�����v����?�dv��oTN֢&@��&�_F�k-��苇��Fe#OOJd֯��|��p��PIQ#�C,0�?��ʉ��%>�rG��M����{����"�2��}��CϾH�)�]�!��	Ǹ�y85�xq���p��F�f�J�2�و_üf�?ǉ�=D�wP�/�w�!�v=��X��/�3/�!X���	�%�% ��5���"�B��2�k�2Mz`��B�@o��[^�}� u��=��5W_~H	��`��,\ަ�It��+g[�N����p$��<
DN͗&8�,�8��!��L�E��w*��ܙw�F�ݚ�Н�rM�e<�!�`�(i3����y�kا0�=<MW�-}�	mp@�s�p���.ᬵy��H��]���ݚ�Н�ss2����
)\Y�����'u���ɿJ��ݚ�Н��W�"�Ů7��B����3�=���!�`�(i3�2*Q=F���q/���<�����7
�e����kn4@Q�/�!�`�(i3k/�z�xEQ���*[UxG!�`�(i3���ꀍ�˺�Q���f�?ǉ�=��9��稕�a�/!O�f�?ǉ�= �@��&}��s�H��rs�i�S�,�>)�_���L����֟DqZo�����2��}���zgm##�^)�G�B�+�WdM4@�&u�)m�$��&;{.�e�<Q���c�ۡ����Ů@�	����W�W}c��ko#��J��Ӊ��@�#��ErS�b�8Z�AԢ�a\��!��a�'�T��~�(��k�C�-�+�g�>U�m��^
/g��6��c�ۡ��sc�̆�!Y����Q�:���Q����.��$���g�e��#����< �R����[�Þ~Q׆��p0̲�2�!���'HY-��
�C�Ʌ��HW�PM�^-q�x�l��1:�N�*�x¥������]n��-��%{.�V#?p�&���A	{K�tU�P!�`�(i3�gCu(o?C!�`�(i3y�Z�;���>0�1ۍ�h �=�f�?ǉ�=��'abW�5�}�]��ϵ��t�pu:�]f�?ǉ�=�O�G?X2���Y �6�ZWq�ߑ|�ݚ�Н��W�"�Ů7�6��,�ݜt���,\ͨ܉p����O,8�ݚ�Н�h�'f R>N0Θ��ݚ�Н�Gظ0����t�%�Z?��<�ry^�%��C����\P�ʊQ:��IK��<[�л���7�~@M��@�Hb�2�Ǐ�t*����B7Ԅ��{k�h�+�0��NZ�Hb�2�Ǐ��t���	�%�% ��5���"�@��A�ی:�Gɩ��I�?g�f&:��r-,l�6>8G���n	l��Q;�im��ȍry��	:��+���������i�����+��cW���}���i����0���LO���){�Ysy�t��P$u��&8�,�oa�}��p�-�o%�'b�be`�t!�`�(i3^P��:w0I� X�1�;LV^Š�r��Lo�_!�`�(i3�2*Q=F�k�mD#V��A��`-2Y��kک�x����y���ݫ�ф���F�)�_�������� "5�]�B�'��a�F�,�U6�Q�L���/��@��:$����z�����	�;�ݚ�Н���"����M몴PBoT�ݚ�Н���_(x��`���^����+�g�>U(��[��`�ݚ�Н�p�n�����^����+�g�>Ub����{��i�X���;_��8W�w��fDp�F�`n��i���-՝-xC�;��|BJ�=$r��H�c�҈��V�ǖ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������;�Ӏ��F�|�^q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڿƿ�d����I����~u����d�}-`e¢Qw�T���P�=���չ���1Y]H]w�
��P��*|u3�M�*A�Ly���Cʬw�S��2����k�k�2y�� <{>w�\��Z�����ZW��<��S����5����.������w���'�(�]�v�<���kv޶Gl��*ң3E�E��'Z*)�?�R��n��h
:h����t�h��W+��W���*�Աߛ+���;aw�4� �ϸ�"^�j���5m��Y�j�`M97��ENҠ����iQ�0�ȷS�J݃��x����Y�iRN���v�Ӿ���yi�1���~!�`�(i3!�`�(i3!�`�(i3Q� ~���.�g3ZrZ�0m�\�O�W,�P �S��n��Ի����\�����ۣz�#˭䱰lM8�!��0�	f$@Dg��5F�*��f�I���s��i	��2��ם� ��u1�|:�i֖��(�^O��C��S�x����6���K����L�4��)�Nc<�tT�!؃H�J�#}�{�~~�^���4�űW��C�G�,Bճ�i��HoQ&�d�k�Si���9��d���f0� ��a`V�.��.�u0��4�ke-t���-���G$��S��n����ěA�E(����h�5,Wlr�r%)cA����L�bB\q��r����>�R�\A��ީ��B��g�W+��W���*�Աߛ+���;aw�4� �ϸ�"^�j���5m��Y�j�`M97��ENҠ����iQ�0�ȷS�J�L�K�vPfÁ��/�6�£wO��l��b}*�ZLN�	���$b4i� ����i9v��խd�g��;�!�`�(i3!�`�(i3!�`�(i3]q>�A�	?�t�ϗ;��|B������kv޶GlR�c4!`��_P��2��@N����(zm�B�q��i�r�Ŏ�]ΟQ��ǺΕR��ӟ-�ЕS�#m,�t��gJB��#U#��F�����p�Q�4���5�O�%E#P[�ɝ�����.V��:��������Y�#Q��~mW3E�-).^QQ���T���b�Bϱ��Z�<��H��h �=��$b4i� ����i9v��խd�g��;�!�`�(i3!�`�(i3!�`�(i3]q>�A�	?�t�ϗ;��|B������kv޶GlR�c4!`��1Z���G&aD�4�X�X�>c�.A�Cw�Hm��p�@OM.IrQ١Ӿ�$pW�q>��97��EN�xÔ_���9j.�l>'�o��&Lt"w��=��Cn��P)�昸�^����yN��7��aq��G�n���t�;���N��I�u7�C䫟۟�>'�o��&L庇�1���m�{��w��p~z�r,7?G)]n�`�I��W�^��D��>�Z�1�!�6��uȪ������:�.�B7�-�6!�`�(i3!�`�(i3!�`�(i3!�`�(i3���l�Nh���W<˥�'ܤ",�����D�-%9*��v�M�{�|L����5m��Y�j�`M4��c�����:/��N��׮	��48ܼ�P���6�5>EZU2��53��(�K�g���yN��7��aq��G�n���t�;���NI	��y7DT?�R��n}�����H�i
�J���̥�0�L�p~z�r,n}_��嗍d&�.�_�L[� �h�����T)#�y�ö�7�-).^QQ#j�o�������԰�W����V'��kd.Cf����)Y����2�g�]@n_���?3B��A���!�`�(i3!�`�(i3!�`�(i3!�`�(i3���l�Nh���W<˥�'ܤ",�����D�-�.}�p'�M�{�|L����5m��Y�j�`M4��c�����:/��N��׮	��48ܼ�P���6�5>EZU2��53��'�פ�G䫟۟�>'�o��&L��)��")�0�=<MW�-}�	mp,��_А#�<om���Ϻ� ��H����8�(�������2*CA>0�1ۍ�h �=���S��B��N�c�B���)%O�lg�;�tb����H�s�
�`�I��W�^��D��>�Z�1�!�MطP�V�n쯎+�ܼ�P����4��Я�g��cH�wA�?ܔnߧ�v;�!�`�(i3!�`�(i3!�`�(i3{�d"����	�,�2Zu����p�����+X��FJ���-&d��]�^���H> �0c���cͧD��_�W�.��;�#��&�qҸ�]b ��)_�32��m�4VGu����p�����+X��FJ���-�g��L*^���H> �0c���cͧD��_�W�.��;�#��&�qҸ�2Mz`���)_�32�`�S��g��I&!y'}��5?�&P-ߕ�L:�,�����^�� !
=�vv�>&KӔ�o�J���" (�P@L0��U�Y��"��5�O�%E#PR��ak����`T�ҩ�	r)��f��X��ͷ(�-�E�u�N����dz����NR�p�'q�-��nEg�N>Z}�C�]��L�溥����v�8:ۛ@W:���#���Fф�Sh�>&KӔ�o�J���" (�P@L0��U�.��/��d�0���.�g3Zꢯ�wv��n�Jt�g���E�*��?�"S���ҩ�	r�/h��c<�+�g�>U�� t��{��X��"��ҩ�	r�_NVT%��y��|Y�
�}I�?d���au | a⣃_B�2Q0��BM�X�X�>M�a���;}`O�k�W&W�f�̒0�.��Y��/z*q+6j�"HsӅ�X��^�Y#ѥh�g8V#��4�|u�eV8���y�)��-aw�n������z��!�`�(i3����;q�M�{�|Lɋ���)���O?������T���b�Bϱ�nQ�rV��q�t7��G��f#��O?���#j�o������6Bj�!�`�(i3!�`�(i3�����z�H{���W�.��A$�P������5d��n4s1�U��B��-";o!��g��Y#&����"sS<�0�zG�������&G�N��W��pp�N1U�)P<�ܓ�Y�������b@����7)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G��+p��qR���Csht��p��Xu���������$��%����ht��p���_���{$f��_Ub��7��G_���;�P�t�5�׹�";o!��g���W�j�T!��w���Pm���֛�l����c�n�RW�A�&hH\� l���E[J��:�����o�.�u:u����<�*%]i�Gφ��<�6�@a� ��fFMqlgd�G}%����3f���K��M�ZP�����Fz��Ԥ�scX{�X!,�'ž1�|�'����u��r��wbk�$`��y+���e��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r��y��j��k��6�
V��͜��!?@K���୩�ݵ�Q�n��T�\ ��� ��g�SE��O�^G�b��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M��ŊPTWo9���=�\;���w�R���yV�'�2\�]��P�),wE�=p��3��P$�Ϙ�O��.��g�]@n_���?3Cy����]E;��|B�]Z#���Ү�6�
V���{_8�Y���d�)bU��O�^G�b��/z*x�n;��|Bs�'��OW'<�w�N������M�U��)���Y;e�iK!���d.���+�^n=\f�5>�.F<!W���t�㮫��r$ɓǃl[�Ƶ�1tSjv�t�R!ME�!�`�(i3!�`�(i3!�`�(i3����;q��b+}y[�6[��u����@~H��k]m��#b|���MJ�a$�Y dN�<@Iv��nt=:��:5A��p&aD�4�X�X�>c�.A�/v�K7%'����;q�{_8�Y��=�}�Vݨ��}Dq�f�v�A�
^^3�V�C��k�HvL)����]�q��I����~uK7͍��|��W&":x��7�֒���dz����NR�p�'q�-��nEg�N>Z�s���Ww���P�|TB��d�hj��m��3��p���H������7Pr��ġ��,�F�����0�5G,��Gc#�����0o� c �ʵ��մHc��,H/���L�����B��2�k1�h�H��*F7	G�<�*��s��ꮂh��,���fR�,� �GR��shbvk~�#x ��M��.ᬵy����uq!\H�q���3��`��R�`�mQ�x�z�oi���:����X�y��s��c�7�wtMM�0�5G,��Gc#�T�Ed!�`�(i3n��>�my$�N��o�/���;7�wtMM�0�5G,��Gc#%@Ԫ�!�`�(i3n��>�my$�N��o�/���;١w��zj�X�X�>M�a���;}`O�k�
�p�	%6n��>�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G��+�t2�G$�ء�!�`�(i3!�`�(i3��}�%DܭOA{�Z.�'�ݚ�Н�&aD�4�X�X�>c�.A��x�`�8�Gl�x����b�'Be�Vj�.�l�x����b�'Be�������H9gUS����a$�/v�A�
^^3�V�C��k�HvL)��+�dr������ɕ�eYl�x����b�'Ben2WȔ�h�U�s
ƺQ׆��p0�Ĝ(�IyI�I�CPWfי�b��}!D̅����<!GO#ݵ�Q�n��T�\ �͉ק��l����@~H��k]m���V'��Kch荛y�(*�6[��u����@~H��k]m����[��N���t/�(�P�/Tu�����_&������n��H&l�x����b�'BeS-�w��H^ܑ��y���8���/��R�E����Q׆��p0�Ĝ(�IyI�h#"�.^��	��uct�td���5N
����\� C&����q��Z��{4++�L�Ѳ�}�%DܭD��_�W�.��;�#s��<�z�0�5G,��Gc#L%BJ�X��b�������Cҷ��ep"�ߏ׍�B��2�k1�h�H��*�1�h�d	�ݚ�Н�u����p�����+X��FJ���-��2n��{q���3��`��R�`K��"���վc7t��B��2�k1�h�H��*L]�f��e���"X��[� ��U,����dz����NR�p�'q�-��n']u4c!�</Sn��/Tu����W`GU�!i&G�\��u������R��ak����`T�ҩ�	r�s�"���A���3A�n�+�sQ}b`�����E���v�RKr�>p�{C��Nq~o@Z�,��#�2
��e�������m[�LEE�S�+�dr����$f��_Ub�F�S�1 �y�}�6f&r#o�]�ʄ�|Nb��'1-/Tu�����_&���iΔ�g�(�l�x����b�'Becc�����4s���.���z'/)�� 0�s],�_�hq`G��Hb�w�2�Q����\}{��E�c���̞���Zt@.���������Gc#0r�϶l���l�%}�Z��1hI����0294l"�[�^��W��kU�%Rd�LCx?�h�����
���PUA�OMM�e�8��
i�c�r׎�m�5h1��0�5G,��Gc#�����0o� c ��4�*ǧ��u��r���#�-�p�@�Af8�ٕ��(�W�!Ċ&���X�G[�T��M�U y����dz����NR�p�'q�-��nEg�N>Z��B|�)�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�s�Yls��8��GM��i��.l�x����b�'Be��/=��v�A�
^^3�V�C��k�HvL)��(o�ܷ������1H}�ɐ��/�Æ��%N����[����2+m��h�����H���ʖ��	�_C*ζ�I����;��P�jcd�LO����K���Yb�Y>�fW�N
%�Rk��4��J^�B^�����f�L��'��UCmV��!jG};�;X�ӛUi]�g�^����H����q���3��`��R�`�mQ�x�z�oi���:��@�����N���!�`�(i3u����p�����+X��FJ���-],��%s��4��D�����C�=�g4�B��2�k1�h�H��*F7	G�<�*z��;S�>������$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx4]�l���׳�D�-p������QQ����"?��A$�P������5d��n4s1�U��B��-Ӫ��*$���A�0rgL�ݦ'ž1�|�'����u��r��m�n���Y�j�`Mx����E2b�z'hۉ)��d�7�q�>�Q�c6�����-ќvlr�{��|e��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����M?��y�!�`�(i3bMGo?� n2ϒ���=��p��N����ȞOߙYĸ-�l[�Ƶ�1tSjv�#2\z��9I��@������˦G�R�c4!`ob.�Y�2W>������$f��_Ub�F�S�1 �-|��Y�$,K�9+�/���p���&Cd�c#��N2D���a{�l�
@\�Zx�.��c�9ʼ��$��:����
�ݚ�Н��>���Dl����|�b�и|��?���a{�w�!]��̍��}Dq�f������!�`�(i3oj�+p�K�J�iN�SE�g�������(ӈ���m�r����fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�Ӫ��*$���A��PN���f;����^F�=�_�7V�o��_�Rv�䩲$��8��I�:Fa�7�����~�Lk݁ 1���tw�i��}�P�|�bs��2[�a��o���H�RtV�^����P%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����M?��y�!�`�(i3����P0����3��x�p�����%>�rGO�D mWN��Ě���aT��3G�IX0F�M;����^FF�Q�f�cny��&���c�IX0F�MV�ҁGG%4vkz����`���φ��<�6�닓.�`�3�P���F\xjzӝ���I(͂��-����q�\E��0�d��+���{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^=@Gp������˃�I�z�iH�Sߜ�*�l8�b(��@��C2K�ǽ$�!b����#�GWW�<om��X|��B�� h�ҩ�?V��j�c��׽���H+�����Dv�/"sB!�`�(i31���~�wӨj]h��J��sr�lE�g�������(ӈ���m�r����fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹���C���NӴ�"�6j�p��b my���=)��r�Ws��(fw���'�̗������k2m�;��|BkCD��9'�u:��_x�'DV���b�z'hۉ)��d�7�qĜ���,�ǰ����adp��e���W�Զ ﭙ]C�1�ɕ7'K[�� ���JH����8����F)�~����H�V�&��<S�G��T8�* � ��IX0F�MV�ҁGG`5:����$�Qu��N.���u!/��"�3ݓ�V�?�f���,(���B�����(�犽{Tɀ��k�V\���"X��[����fbK7͍��|��W&":cp6Dq��;���EWr�4br���Y$�J��;xZ��j�
�iB{�Z�_��?� Zh�R?�R��n��am�Za(􆿳��$�Y� ��l|�*"k���(ӈ���m�r�����$�Qu�9s� l�XF;p�	_�S�
utY�{'%s��jb�ܳ���p��b���a�'U^\�T�\ �͓D+���4YV����(K7͍��|��W&":������y�:Fa�7�����~�Lk݁ 1���tw�i��scX{�X!,�'ž1�|�'����u��r��V�ؗ�X`u!/��"-[���V~e��0�U+�qbp@�!�`�(i3�4br���Y$�J��;�ˇ�h��<�W�.�P�	��
�Q�}hs�����F;p�	��0FB$��e��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r���'��o�u:��_x�|�\V��]�!��	Ǹ�y85��iV�����~�F�
�ݚ�Н�|�au�(ZԵD��0�r������ҭu:��_xBrsjUd��!�`�(i36��J��c��Yu��^��.�mZ����w�z�'�P��yN��7��aq��zW�&��F�u��r��!�`�(i3���e�T�%�td7��͝����ک��l�K�>�������Ra])n#��Nh�=f[��8��GM?��.��U��@�fћWQ�g��	�0�=<MW�-}�	mp5���%�+� h�ҩι�+�t2��&����!����omi7xK7͍��|��W&":�ݚ�Н��H�����4br���W��Š��Օ��qvdЧ^{�jMdGN���!�`�(i3�'��o�P�nq�S���i
�P�nq�S��%���!�`�(i3��w�w:�!�`�(i3�'��o�P�nq�S�/�O�Ha��my$�N��o�/���;!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx?�@� !D7Y'��k�r�Ua�;��|B��loXB�R�S��>j���(�'�'���F�