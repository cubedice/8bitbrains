��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	��q5.A��|�H����VM.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I+ĂiW,���D�+y_�L_H��-..i=?�m��+�<4��ˌ��|��v��ӳ��$Fe@���N�w	*D���y&�f��+K��[y��ڂb�nP	�'~�e�r:���/lt�3� P�;��1�-���/�_m��37tw�n�&/uP!ߌ��˼�{�&�z(ݲm@�)yH�I@'�ew2�\�蝆�u����l�|���j����1�}�<RK��2Ee�Y�R2
�I.��	���
�Ɛ��BR�[_i����v H�$�Yo�1z�:맷�m��d�78�^f��G�n�QX�v����<.���+��T���jB�Fg�:S�Q�[�$A�������6��H4�
� �AH�T�t��3��'�Wا[~�l]ǜ�����] ��F@�4%���D�Pfc����2P����/�"��< ���X�M+��tc��P9P��`�.�D���J7"�x�YW��t��⫓���RL�a)�O��u����H7�Q?�"�B�gf|��q�7C��H���j�v�?�r	⚎���k�8���҆�|n���u� �(���.C����yY��:J�Й�m��C��ߊk'�4+.���`uI�[l٧cJ�^j�u��w)�S��X3���7��Mv�9�<��{�d	�I�
y�8�:r&@�bD�	)��m�D=V��R��c�ȸ���T�٥��T�Sҥ��|E�EYZ/�J�|(��jrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�T�`�7?�ex�`����gZl�B��E�Wm�g�X��ˆk�=���;�w�ln'!MXi9�
���s��3{�β��CE<S�In'�J�gy�	���q�Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S�7���I䟹�%H�$��ī�o��<�)�G!�u�����!�M��EE$ô&y�uZoO�=���@$"��ea�8���*���g S�7���I�t,:=g�B3����Ӥm��+���uN�YW	��V �T�QT�8���v���I�Uu��i����*�{¥������z�)
ԏ�.T٢ߡ[p40�zɈ:��B��J��H9'E�HG.���hm�F!�`�(i3���P!�&K�A�H����8DE��	�J�ILo�����,[$�	J���GKer�I�F�ݦh�z�(������l#��䩛���y��lD&خ.�o�O
��^O��w��ԩ9����'*D�]:�W�G����?+D���0�7a
��r�yد�9�����~���-�f�t�������~��(,R[#�(y�T%ME)��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3o�kr�.z�o��x�v!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=ؿ�?��5Q�Ub���Ɩ���2�Q��0m �]vo/~�e6j���-M+�Ԝ�}Dq�f�!�`�(i3!�`�(i3!�`�(i3!�`�(i3zZk���?,�=k���52p�8s�?�������`F�k�d�l�!�`�(i3!�`�(i3!�`�(i3!�`�(i3(2��\YV6{,q3�+���C��n*�k`��ͯ�K����6��~�?Q!�`�(i3!�`�(i3!�`�(i3!�`�(i3_Q1������t?uw|`�ڛ�m��e����2��=!�������Mڂ+!�`�(i3!�`�(i3!�`�(i3!�`�(i3�1�?	/�V�8��/��6�?��h�0�����9��S]��ݚ�Н�:��9KmR�^Ƒ�Ӈ��t�9>yh��DvO���v"�N-�T�\3%/��.�@��RN�]�5'c`�/��ȍry��	�s�٩�삠k�bWbG@���p���ݚ�Н���?��[� �V8��v ʞ���
�:qEp� LTx%�0�أ�Mft�s� u�?D�8�镁�aR�!�`�(i3�i����u��N�v{���df"�	-7���C��L�c27���&�_��lC��U7�C��zC@��f��p�(p���	��
�Q�}"�4��m�S⏸[��]2�y��]�!��	Ǹ�y85��9�L�fG"j���b7Z�n��[��{_8�Y��=�}�Vݨ��}Dq�f�i�]ʺ�
ǳ��ٜ�]Ǧ�JS�cbp��'@
9��y��5�%]�����3�(���tP"7��%e��0�UX�Pp42JF��c;x�@Ã�D譸3L�*}F�x�����Z鎬����Ĺ#{����}Dq�f�)�{6�U���ea��L��K�*� ���G1��[��K�+EC�����6��lC��U7�C��zC@��f��p�(p���	��
�Q�}�d4�n�Yct_��צ��
t��{<���낌)P<�ܓ�Y���aR�!�`�(i3m����'K���Æ6�HaDl��+BY��9��8������{r��;�¬pX����B����qe�@Rv���|z�ä�@��m�r�����I���`��`�v����2y��l����4�n���xǊ�Jם��t&:���a��2��1�V����(��8fDs;ly��\%��'T���+��^�Y_Ez��!%���Kv���ft�s� uƍ2���lğMg$9�rJ
_�y�V( �w�;>cbp��'�����C��ݚ�Н��l��#�}��
�'����j��<ͧ�:|��b+}y[���S�fDV��,�����
�9�j���B]��>��y���|e"�7؛ڇ��lԇ�-{�(��̓i��:|[%.�|Tck�=�mJ�0�6��q�1Ig�I�?g�f�(�r���`�s��;#�A�v��
~�d���	OQ���.rA�q"�#�)ޒ1�:�Ω�q��� �����_N���m3��>�@�;`)�;�$�&��[�@*`s8�R�	��_X�[��l����4_&���&5�(1Lô �ԟ���7�����uhP��9�j���B�<Vo�eo���9�r7�K6�L+�.8ޭ�;���E�qA��~��.�f�n�f�9�j���B0���\,�2tW鳲��u)+�*���o�7� ʞ����H� }��|UY/
9D]2σܕ�4J&)��͈H��<d�x� �q#�W��=A��$��mNw'L$�����/W�1�䉁 �?,MU���k]m�����i�#Ѻ'���Xw�j�7���+[��@yc�&ck���CyW�f�t��ł�!r�dN�<@Iv��nt=:�i3�|)sՀg�u�+��yۂ�J1���i�#Ѻ'���Xw�j�7���5�%]���a(􆿳�tP"7��%e��0�U+�qbp@��dט�w��l�,�9P��Jw�TI�~P�b`�6�Ƌ��X���`��w�K�ʌ���p5�]���7'�o�$C�|�6soi���{r�����ތ�1ʆ�In��t�\aьIR=Ϊ�/-T��G㏐���g�,P�n�U���q�
@�<[n^/���\�e�$�L� s�j8�҇D��μz��z�������f�62�-�x�k��V�4����,D<���h]��/�8Pxκ�ǣS�\�m���k��V�4��)�,5���A\�5H��߷~��nJ!-��|'U$I����A{�c�!5�k�d=��¾ȼ`�����t}�T$"��ð��T��vr���I����}�N�<�>��LҒ �ѝ�:���y��lD���	ĭ<�����Km�F�1�I߾��ٸ�(�!�`�(i3��Պm��%�1$��ED�2�Q���K�V�!�`�(i3<.�cs����!~f�{�e��@�	m�Im��/9�=eF�ѳ��{|�B�A��Z���Ӗ�����G�k9[b;�J_w"�7sG��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3cW���%�	t��C'�ʁ�;C��l6�P��{�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л���O�/=1�u\2[�rNj�7��9���r����!�`�(i3!�`�(i3!�`�(i3!�`�(i3Y�4Eb�����@��G�ϧr&�8�] ba�Mg�wì^�3�%�X�*�I�����o���ڻC�i�φ��<�6��֍z����!@�Y��t�|�AS��U��)���2#z�Ľz�`f���sd=��¾ȼ-�,A��g�ΰ-��3���-����!�`�(i3g�F�W�k	䶙%���K͸�6K��7l,%�z�-uͺʉK�/�n�r���pu͟0S��ϐ�LD��B�r�ve/��I�3,l5�wK��&�@�	���Ĕ׹��L<C%`�P�����
xM�v.����V�8�|u6���H��y�ћ����iH�}�g�"{��n����8-|�DU�
{�~j4��ۊ`fSc�o$NG�&ց�*�i����D�ݚ�Н�B�%@;V�䜯}Dq�f���dEߦ���m:���q9+t�}�ݚ�Н��k��M�RK�a��R#	�N�QT��a��o���H�RtV�^
��X��F��[�i�[,CLЈ��՝� s�#���k$ ��+D��HBڎ@L��LT��]
�:qEp�;�P�t�5ʁ���Mյ��Xf6�h��ݚ�Н��{}yN���?D�8��Mg$9�r;��`�x�����6N�ƺ'���g��+��9,(bulx���a��o���H�RtV�^
��X���W��Pw-w���nNH!�`�(i31���~��'T���+�N_��ʥ���Y� �����"�$f��_Ub����pT����'��@�my$�N��ݚ�Н�6Gި���74/���
8�	3�����1��ݘ����$�)�vx�/���)�G�rA���r5��g��(�IX0F�MFtU�'�!�b_�HN�d
z��n=\f�5>�OV�vG�[ƛ?�	�y��xZ�&J�:_7�O�����WS�;���>e-Gb��F�%��v��`
 ֢���V�ܔ�s
�����z�+��9,(�P�U��k��-����P#+_]ݱ��3,l5�k	䶙%A��ʺ�l�������B�'��a�]l�B�:	74/���~:�*�$f��_Ub��}(���603�gea\�3��Y$���ܡJ��0'�^����/�"����y?�Yam�"�"��ӌ�r`���*1i#\��u��.d�i�>1tSjv�c�@���Pxκ�ǣ���Y� �����"���jVѭ@P#+_]ݱ��3,l5�k	䶙%�F�}қ~���Ě���M��%�p@t�td���5� ��F���}ō�X�]l�B�:	74/���
8�	3�AL(�z��QΰU�P!2�͞nOY4Px^̝�_���s	 ju�0�T���A��!�|'U$I����A{�c�!5�k���èV����94��؛1tSjv�J-ڦ�.�5��R&��dN�<@Iv��nt=:�oR��mԶ�4 >y�;o�� ����nF���<�W�.�P�9�4��ow+\v'�]5ʈy�@�oI�(�w�Q�� #�	�';��#j�7�癆cg��߹9$���9s�{�����&G�I���`�v1a{J��;�Hf�MN*�����������4 >y�;o�� ��'*�ha�u?��F�zw�}�	76�&�� Ӗ�t�c,�\���$�)�vx��=�)�r_���s	 j��̇��'_���s	 jR2,#�����`�v�˳V�0Kg�:#�R_����J�����m�XQ��À��`񚷱��`�v��"��gL
ETk/�0�������f4T߅4&b�ՓG6|=TElJ�̆% ��J��ɞ}�UBW��ɯ��[�҃]U���Hr��2�?F~4�0�*��� �B�؜"�37�˱�5�7F��%�%ح�e!d�\4x��'k��l�����{��\�'8�쐩�8toC1�Yܕ~���kR$��h����k�xU����_�8���< @���-��00��;ӫ�j�5��mz�0�(,�FM��L�Ex�e�R\�����S��Bb+����6eG����V�����a�D2Z�+o9�t�Wm^� �L^�xv!���wH͔I�=�=F���ˏ��Z���+]���P��@��~h�{_8�Y���˂lq��qgF���~Cy;"-���!O��ʅ�UE�TLP
���V�,�=R�/���H�V������R���YƼ/sf�e�}s�dKa���c��,�)$�v1a{J����n�#+=�{r��;�¬pX��g��U-�e�wpb�Q�`�|��K�z>���@]����ٲ@	�*q*�K?�d���&��ǣ�W?����4(/W+�����ڻ$�춵Q17�b�����d���!iB�6o�ə��:X���my$�N��+ �Ę]V��	��y��J��[���D������Fy�׉��
d�YB%��Wf��K�;��|B <�Az��'\��i�J-ڦ�.�5ɠD(c!)`�|��K�z�5�%]���a(􆿳�f�(�<c@;��|Bz�$6���{�]c�h�ʔir��#j�MJ�=��7