��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�"� r��������:N<��;���Z��4d��{�
��|��Ȋ)zo1���á-�w~��d�������mo�����(����5�a���V��$.:&R�nU���T���딣0&_���X0���2|	p��rw@	@us���)�]&��_	��u|��yq�`݊�|���"rG�
���}�\�bJ(9�{��r�H�����طǪh��p��U>?���>�`\��Yi���u����l�|���j@��"�O��$� ���xI+r�� 0�D�A�f�mXׂ�(ѳsv�`�S��Y�ix�P�Ra����+��a̞w���{ֱ@�W�8d4؇��2O��'HY-����T-Q3�Y�h��~�a��9�ĒTC��0���Gʺ��7F_�X���h�W9��U��b��j�\�����OU險"Ya��Aq�[K[n�8�����F�H�h����op!!v*!��ċ�G�iNqϕ/67��b"����S+0sY��<�.�zn�"Cݪi0i�����V�YB�H��ٳ�Xݣ�(��Œ5J�2_[�!	�^��ܶ2�s��b��<�vd�̪��g�}s��4dr�)w��6�J}�	�$F5�����i�-
T�����N���RU���	x]�<��O~��z,}�K;�38��ɓE��m���>Ly��V8�-P����6rG��>zX6AE�v�hH,`���s��8	R�s�$tA���]T���ɨVu��7���	x]�/�Roȕ=�~篟|�nNMR�ȷF��θX(�aa�y����g
aC��eb��T�Q5�Mt.K8��~�X,.:8GT���1�w�Ҕm����G}�ھ>�g��u��w)�S����w�~篟|��1�`ߘ��J�P�aa�y����g
aC��eb��T�Q5fs7%=H�n��>v����u���Lo������%���]��\�4�sP	�b\qB�xy�V�2yE�W��rE�]7t۸�~�MUs �.Eٓ�9PHvE�	�����}�m�!=�y����h�}�{Sh�xy�V��ԋ���w�E��"�̣��}\l���?ڛ^T�k��e���p�c�TQ١Ӿ�$�^go���y���2���=���'0�k�8���҆�|n��5����s�!���3�@�VIg��5#���H	��Ŀ� [U ����k�ә�3-v��Q%RH�,�@&�Z~�a�0�ߋH������<
u��������;1��
:0�[�H^�*K��$�U���=��-]d�yv`�m�����r�O��C��0���[�	�P���I�W3V��#ɐV����{D�\�����e0���0�YՕ�j&�S�i��G��RL�a)8��Q̮�D�-��]�"��3�����;H����U��Pa�i��TH��O��R��c�č���@�,�AQ�CE��0�̀*� :��������|����`��h˚.��U����X�U?��f?��w(�]�k�8���҆�|n���f�S�z�����FT��vY�]e�u�z��[�_yǨ�7&s�7�L����ݲ]�mCu��w)�S��X3���p9�AE���?��|:0�4��:uD��B��z�J�d{��Z)C� Qܤ#֭����RL�a)8��Q̮�F�������~��j�n�?��;H����`�ü
�*�`��#B���l�t��m�!=�y����h�}��a_qz�8Y�&�\��-�f�M��	8�.)��hbHp|��Û���_�:Y���k�8���҆�|n���:�o�E��Uu-M�rt�d{��}lJ�Й�m��?�Vޱ������{����VjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�׍E�+��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E/?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_E$ô&y�����[�/�H*�m��/2�ޅ���?�y��h��ؒ3����]ͧF���y: �����v'gn�]o��in�m��+������R$��Ct�z&��ÃlO ܅d��
�b�lr�r%)cA�����Y%T��BP��&��J�'����IEߺW�L�sQd�h�=3�!�`�(i3�i3<�f�D���X���`��������I7��-5�B�wj$g!�`�(i3�a�\����9�	��%
a���+P��_,��ޯ#Q �4�M�����jݭ�F���L�D��6S��X�u��
)\Y��!�`�(i3�E����F���8�TP��Vchw�D��y.y�Q\�@vs""��Fq/�bi��±�sR�{F3�_� ������,��\G�Y?�� ��}r�x�e�X�����5	���]���c�A�L'��!�a��5�%]���a(􆿳����^��$���]׽������E��@IE�U����S8�/ #O�)R�^Ƒ����"X��[��Q[R�7��=m緒��J���W�7G#+�Ǘ0z�cULd�g>57<�C�u)�6�3A�)OqЈ�&��g3�g��U-�e�,���6+�_������"B��$I��w��,c�A�L'Qī�*pY��㶢�&-���x�'@�(��P�G�p�P�į�d��8���/������T!�G���-N�By3��<�]�!����M[��Ǣ ��$�,�������5	���]���>����C�*��^�"~H7.�;AF@IE�U��>��l%i�-]a%ڔ��E����F7G#+��\w��0]C$mQ��"�,�>E����-��%Mό���.��_F�k-�!�`�(i3c��Et��q���U�ЂDa��(o��0��7��|g�Y�'���Xw�E�i�m}6	��	Mk�rv�ј�"��Z鎬����y��|�!�p�tN2s���(����5�a���V����L��]�>}|��XH�����,>$+W��� j�(����5�a���V������h+=:j�r��VYW\��+�y�^v�㸒8Kq�b9�����9B7��Q!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����Bg涆7���ө�)�F��3A�)Oq�fhz�����bu!�G�Ḁ� >e��{�,����*�X,JHn��z��x�f7﹏!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3͈�
�b�̞��>��bTg�zϾ7���q�>�$��Xo��&<ՎL��W&�C��.��lJ��튝�b�Bϱ���w�K����+��dЧ^{�j$��XCp=8�b(��;3��o�r��Cҷ��e+�6��? �B�P��w(��7���ө�)�F��3A�)Oq���(���B��ɓ�~Ҡ	��[�)�D#���ߔk�V\�V�֓X	�@����gG�?#dK1"Sr��3��ő��̼xZ��j�
�iB{�Z�_��?� Zh�RG�p�PR��{�&�8���/����,D$ů6j�e���;��U�� ��q��T�ٮ|�,
����$C�~x���yM��?IK��y�8���/�I����"�*�şxˏ15K�@�/�d�٣��c�A�L'Qī�*pY��?� Zh�RG�p�P�"i<,��1��yM�׶��	��:�g��U-�e,%�0g���j�|�{'�XYS��q��T�ٮ|�,
���A�;�֋`N��7�j2��'Kb�|n���7���ө�O6�]Η^a(􆿳���2����.〧I����@�k��}�U,�(�)8���0y�	�C�u)�6�3A�)Oq�fhz���I�Ūeߋ٣�o{�i7�v�ԯ��Q[R�7d�x� �q:��j�g��$�K��{Z��rs�i���`�M�	=̞��>���ԜF�����`���W�L�sQ������f���[��R|#9���b!��u፯����n����ȼ����f���,(���B���ި�����|`��'��>�4Nu{ᵿ����-R�4���d�a�4$�b!��u�;+�'ն������q��T����<�սѡ��`y����@����gG�����5_�6���9(�UtW�*XF&|S���T�\ ������q�f@�pH�:V�^3rdS��"�,�>E���]�!����w�Հ�b02�OQzg� ���"�,�>E���]�!����w�Հ㋚!iW=�!�`�(i3"�,�>E���]�!����w�Հ��zly�Ղ�zM#��m�"�,�>E���]�!����w�Հ��p�04�/���jP4J�"�,�>E���]�!����w�Հ�[�=�5x��_�Sc��"�,�>E���]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e,%�0g���[�=�5x���_�*8�"�,�>E���]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e,%�0g���[�=�5x�����c�"�,�>E���]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e,%�0g����ʐ��$���Z��owGT��p��]�!��	Ǹ�y85�B���0���^̽1��R��ӟ-�F`���G���`y���!9q�OA�^V#��i�9�/RsvL�!�`�(i3�����,��(uB��m��I���6k��{��`���HW4�wvA�qS�F_���ٱ'W�w��fD묈�϶H6�9Ae L�x�S~p�A�W/��Wu���t�T��?E-h��$^(?��"��h��w���`���φ��<�6��Lt���hm�(��k8��ʡ.>�xjzӝ���I(͂�'�ɳ��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g!�`�(i3�����n��)��RU��my$�N�����X8�՝� s�#0�ʂ�j�Ï��	�l�lM�3 zM#��m�.�
9� ���(ٗ.;���JTv���H����o�γ�ha��o���H�RtV�^��#�a�Ą1 �u�.������&G!�`�(i3Q3S����,1��m��xx����E2b�z'hۉ)��d�7�q�!�`�(i31���~!�`�(i3�y�3�����$PW~.!�`�(i3�G'�a@�{~1JS�K{ð��T�ݚ�Н�����l��A·�a���ڌ�&-���x�'@�(��P�G�p�Pۙ�Wl��pH�RtV�^!�`�(i397*�SCu̀A�pi�x�q������'�F������!�`�(i3$f��_Ub�F�S�1 �
�:qEp�;�P�t�5!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;���⾰��J;_Q���Q�X�G[�r�J~��ɥV��	��yq(��q���J!�U�e�v2�l[��Ģ�e9Y��s7"�,�>E���H!��\s�(uB��m��I���6k��{��`���HW4�wvA�qS�F_���ٱ'W�w��fDg2K��O����,�����n��
/��y;��`2����]'\gWg��	�Z�kfc��2���8���+�^n=\f�5>���1ë�LA��R�ߋX8%�v&2\���F�`yx�>�+X�[�G���K!�`�(i3<�6�Q=��S<����K��!L��3w #�T�Z��&�2����97*�SCu̀A�pK7͍��|��W&":VA�ڦ�c4����g�Z��3��a���!@�f")z.��W�����F�P�7��S��h��d\�����l����� �'����u��r��;�jmT�#Q���V�_�mS8<�n�ݚ�Н��Կ���p5��6V�|��nF���<�W�.�P�	��
�Q�}՝� s�#�=����T!�`�(i3���ifz�d=+ӓ��#!�`�(i3>����a�����%�g!���2�(!�S_�gWaU �IH�RtV�^!�`�(i3*��0st�7�j��B!�`�(i3��i��:q�5/�V�q2P`��� Z�y��	�����u��r��!�`�(i3*�˜	����r"nCo��I�Ūe�ǩ"�4s2��ԜF��v��?���(�
nЯ�O�!�`�(i3H\wN+����&$?���I�Ūe�ǩ"�4s2��ԜF��v��?���(�
nЯ�O�!�`�(i3H\wN+���S=��-��I�Ūe�ǩ"�4s2��ԜF��v��?���(�
nЯ�O�!�`�(i3���v²*^�:�6�'�K1Y�q��؇�M.9j�֎���x��y�o�!�`�(i3!�`�(i3�����n�����h�&m����fJ�1D1�_'���p>�!�!�`�(i3���%>�rGO�D mWN!�`�(i3�k��^�1��������u�t���Y�;���U;S����xQ�1tSjv�!�`�(i3Q3S����,1��m��xq��c�3�+���F��ݚ�Н��Ra])n#���r����!�`�(i3��^x��A'��]�ꛣ��yM�B(p`D҉̖�7�j2�٨%��W� ��ݚ�Н�!�`�(i3-����p�ȐhJτRgR��yM�B(p`D҉̖�7�j2�٨%��W� ��ݚ�Н�!�`�(i3-����p�ȟ&�h��g]��yM�B(p`D҉̖�7�j2�٨%��W� ��ݚ�Н�!�`�(i3�rag�S�m������4�uJ3Mu��^3rdS����4y��ij��-����!�`�(i3?�k�V�?����fJ�r{�-� ��]�(ld5��(<��e؎��z+
!�`�(i3���%>�rGO�D mWN!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ�c^����24���7�T�O�.�g3Z�)V��B�1���k�}�����iso��8���SY�N�W/��Wu]���o�)6�o8:4�I���c�90�Ǘa��x���+�^n=\f�5>�܇1~�}��Eg�N>Z�C��$]KC���"sS<�0�zG����ZAL�:!�`�(i3���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+�#}�{�@�m�W#��H��97��EN�Q,�SGŹ�R���Z�F�\Ȳ�r�r%)cA�n��If���8�6�e���;��U�� ���^E4+у��b�Bϱ��MQ�'����㶢�&-���xԲ�Z��*����Mڷ�2v.^࣡N!�`�(i3iŞ�W�%3AԢ�a\�ɓ�~Ҡ	6d�dG�7:�R���Z�F�\Ȳ�r�r%)cA�%�\B�����x.�KnqQ�����(�6k�4d�-��(�Ļ4��aA�'�I����~u!�>!��N
������U�� ��!�`�(i3� ��U�_:�>=:9_�ak+Q�h'�Ȝx�5W ��̫(�8�u?��I���?B��#Ɵe�*|�÷�Wе ;�jmT�#��"����G��Hb� h�ҩΏ��^Kho�7�j�Γ��-����!�`�(i3�kv޶Gl�e���;���
`_�{_8�Y��=�}�Vݨ��}Dq�f�H�5Bj��@�m�W#��.P5�iŞ�W�%3AԢ�a\�ӄw����$C�~x���yM�we��k�)!�`�(i3K�\7}�W,б �A	�J�a$�Y 97��EN�y�JB���P��7�j2�ف������̞��>���ԜF�����`���W�L�sQ������f�E��3!�`�(i3Y[�Yy�l�Y�F��(�����;qn�)�� �g!�`�(i3�\d:0�g��
z�.�MJ�a$�Y ״$(�>g�
�:qEp����p俚��+�t2��Zh|����q9+t�}�ݚ�Н��$VǽO����D�D�����r����\���F�`yL��.1M?��y��ݚ�Н��H����� ʋ�aGM�о٫��x>O� &-���xԾ�J��RQH�RtV�^!�`�(i3� ʋ�aGM�о٫��m���\�n�my$�N��o�/���;!�`�(i3��w�w:�!�`�(i3,\ͨ܉p�u-/���y�8��C"���o�k��e�@�m�W#�:gLFX?�]��}Dq�f����%>�rG�@�	����!�`�(i3�3�7d`yu-/���y�8��C"��cG���`ö8�b(��MdGN���!�`�(i3;�jmT�#�#}�{�@�m�W#�UK���6����>�4No)�T*�c���-/a8!�`�(i3�B�'��a���p��b���ez8�US������`�K7͍��|��W&":�ݚ�Н�
�:qEp'{w#/ B!�`�(i3hs�����F;p�	+��Q��:~fz��ro�)���Z��oGM�о٫�1M�.(*��!�`�(i3HN��R��bP�63Z�t!�`�(i3�5ߧE4���ݚ�Н��H����� ʋ�aGM�о٫��x>O� &-���xԾ�J��RQH�RtV�^!�`�(i3�⵽2�RH<�2�8��C"���\hw�h��r�r%)cA/�r�]/2�ݚ�Н�!�`�(i3��۵��(2v.^࣡N��4FF����w�FB��-/a8!�`�(i3!�`�(i3K�\7}�W,б �A	�x����E2b�z'hۉ)��d�7�q�!�`�(i3!�`�(i3Y[�Yy�l�Y�F��(��įէ3��}Dq�f�!�`�(i3�����!�`�(i3!�`�(i3K�\7}�W,б �A	��s���6�XYS��6 y2��R�!�`�(i3�y��j��k�����5����j�)��ȭzB��6���91M�.(*��!�`�(i3���%>�rG�@�	����!�`�(i3�Ra])n#���r����!�`�(i3�⒍~���yp[ E$�K�\7}�W,{�2|+wh��7���ө��.Y��(��ԜF��g.�~R�>������!�`�(i3���F��O��ݚ�Н��Ra])n#���r����!�`�(i3�5?�&P-���P�/�cK�\7}�W,�b1��G�p�P���� �!�`�(i3���F��O��ݚ�Н�$f��_Ub����pT�HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}Ĳ�y��iE��ez8�US������V}���]�p��Eg�N>Z�`2����]'\gWg��	�Z�kfc�?)zni��`���φ��<�6���')��8#�W/��Wu�7�癆cgQw�c4~Nr_�mS8<�n!�`�(i3!�`�(i3}�gv�oE�[��s�A>�xw'��M�v�����FK��|�H��4"�$�`V1���j;9ekE�g�������(ӈ���m�r�������F1��h��;��įէ3��}Dq�f������A%=�Bt�^�>d�g�K�̢k���F�KD�Vr[/}>5��0�7<(�lb����y��lD�7m�T��Ʈ+ˀa��z��2�,�$XR�QܛOcOZail������&G����l��P��n�#�$a��o���H�RtV�^9��?xs���}�ڍ�����;q�{_8�Y��=�}�Vݨ��}Dq�f�a3@��[/���fg�p5�+�}�OGn�)�� �g!�`�(i3�>�u��8f��P����k���������|e"��w�w:�!�`�(i3�c��;C �3<M!�`�(i3,&���	�)��ҕ1�PS��-����!�`�(i3�k'��e�ؕ�22�� ��U�_:��}Dq�f�;�jmT�#���D)��{��G���ϗ�\��MdGN���!�`�(i3`
 ֢���@�k��}/ ���we��0�U+�qbp@�!�`�(i3�	��x��ݚ�Н���6�����7*9uu�I����~u̲�2�!�����M�!�`�(i3���F��O��ݚ�Н��H����̲�2�!�P����p��ݚ�Н���6����Αk�]I���,��~!�>!��!�`�(i3�k��^�1̲�2�!ڄ�]���J���S�<Ԣ�7Z�:1�\mdЧ^{�j��-����!�`�(i3a3@��[/���fg�p5�
�	��� ��8���&�
�:qEp�h?�4DM3-���~�$��XCp=8�b(���sjߢiVr�r%)cA9��9dJ�!�`�(i3���Ȋ�?Ӗ	W��e��*}�T�z�D�R!�`�(i3^��4�Ј��r"nCo�o��h��x.�Knqd��^��R��ӟ-�%�ɍ��=!�`�(i3`
 ֢��.��� j�H]���ݼ�X8e��e!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vxgd�a�"�
�X�G[����O��6O���N�S`��ޥ��IX0F�MV�ҁGG�.Mm-;�d�G}%����3flLnN1(�ZR���:���^��@��'ž1�|�'����z.��W��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g}�;��������/s9����;q�"��ӌ�rɎ�#���?\a��4諞ic)�̩ƍ2���l�����g�Z��3��a���!@�f")z.��W����Q�Y�;y��v��\���
^�|#HK������ �'����u��r����#�a�Ą1 �u�.������&G!�`�(i3��JתMܥ�I����~u���NM�����'T���+��PJU����-a0a3����|e"��w�w:��ݚ�Н��G'�a@���Αk�]I��w��FR�-��(�Ļ�ۈ��ae�O���Z>m.��� eoK�UuA�����5����;��ɻ҂�V�'�M���V��+��Q��:~����t�Ƥ�x.�Knql5R?}�b��2��G�Sr��3��ő��̼(�̖edЧ^{�j�ag:zdu�����P�<z'�$쾹KK���������E�§"�p��~u��r��!�`�(i3�G����ic)�̩�?D�8��՝� s�#���k$ 
�:qEp0���Y$�k���������|e"fĉ>99��A0ok�ª���l��U�����9�;�-mO��ȭzB��6���9Ns�ﭝ�H�RtV�^�F{/�����,([�y���8.��휯}Dq�f��	��x��ݚ�Н��*������Э~���V�q9+t�}�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx+���B��d5%����8�G.`����).�
�]�!��	Ǹ�y85�}q��m�l���9�b:m�X`�7���ө�)�F��3A�)Oqn�����ea�g��U-�eFR��9�o��$ BŊ���/x�c�_B)+��=����Q{s�	�R��~�[o����D6�~�ݵ|��*뇺�ѯ���Z¿i!��j9�7�awf�{�p��ν(C�.��[�}�s�扃�+�z�.��"�]'\gWg��	�Z�kfc�?)zni��`���φ��<�6�s�扃�+����F�	A(�c���_G��Hb�8�u?��I!�`�(i3�d���a؅q$��.��m�f.���G�?v��� �+��R��?V��j�c�_�Sc���I����~uK7͍��|��W&":����@|����^a�nu4Bޗ��jw�	��!�`�(i3lG%��`��ǚ��ظ
��@�U#�s�Yls�<Ԍj��_�mS8<�n�ݚ�Н������y��'����u��r���2��}���4�a1&sx����E2b�z'hۉ)��d�7�q�՝� s�#���k$ �H����/N2~-ٲ�5��X1tSjv�!�`�(i3�)���IrmP���v�}�b�Ot�i.�\��$�fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�����A�;�ˡ��>O<f��J�'8��dA�IX0F�MV�ҁGG�.Mm-;�d�G}%����3f���K��M�#�Ycм5����"sS<�0�zG����ZAL�:!�`�(i3���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+�#}�{��Y$�J��;!�`�(i3E�g�������(ӈ���m�r����|�au�(Z�!��w��v�~/��n��>�my$�N��o�/���;��0���>����jP4J�!�`�(i3�I����~u/��kOT*qA����6\�4�@�� �-jېI�q������ л��E�BS�+��U�,�P!6���r����L�J)���� \L�1tSjv��H�������bO��M?��y�!�`�(i3��=m緒�6�T5.Ze����;q�{_8�Y��=�}�Vݨ��}Dq�f�hs�����F;p�	��Œ��S��nF���<�W�.�P�	��
�Q�}</Sn����+hX~!�`�(i3��$�\%e��}Dq�f������!�`�(i3�#}�{��Y$�J��;�I����~u�kv޶Gl���m\g.�\��$��H����5/�V�q2_�mS8<�n�ݚ�Н���(1l�jG���Z��o�Ry�����!���c�A�L')�_��rH<�2�8��C"���:5A��pfĉ>99��A0ok�/��@���@!�mg?!�`�(i3^�R���c첖�7�H)fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�����A�;��e���Ԏ
m�S�t��K!�`�(i3'�^����7>`[�J�a$�Y ^���H> ��n�U|��%�-�C��7�Y &����"�`y4k���Z!���C�H�>G�g������1@z���rs�i��w��V�H�N,��⒍~���~�]���]�!��	Ǹ�y85���?�A��	����wN+�w�2��|F����y
���S���F�,�֏��9�GͿK����S���� "5�]SƏw0���D ML:�,�Xʚ@h!�`�(i3!�`�(i3fC��T����ܼ�s�٩���I���Т��^�\!�`�(i3-��qW8+���ǣ©��qr�^*4y-��u)+�*6�X�$�!�`�(i3���K�7���[�쮃���=����t��cg3/F�~f���|�H.z!�`�(i3�b[�u2�Gp��bە��Y��j3��� Q�N��*�������,�Xʚ@h!�`�(i3,��O^�{	��O� m5��@�hGq6��nX��U�	vn�����7Z��-��������o��?ʢ��r����`�4,�pI�!�`�(i3!�`�(i3!�`�(i3��g��E��� ����N�v*$�!�`�(i3!�`�(i3!�`�(i3�f8Y><&��\��f�?ǉ�=���gRI/,�Xʚ@h!�`�(i3!�`�(i3���Z�N�j����t���hQ�GvE�|43��52נ޼��X�B��+ H!�`�(i3-��UR5�(<�%by&6����!s�;�����,�Xʚ@h!�`�(i3�&8�,���rRV��E���ci���Wʁ�w�*�fBg�!�`�(i3!�`�(i3�X;p`�FJ���f�?ǉ�=!��I\+��M�a5��|���瀆!�`�(i3��L	�����T-�l�����b���V�Lx{<qH�~�!�`�(i3!�`�(i3fC��T����ܼ�SSB�����m�%��~?H�?���i�jw�j���[��c0�]�:�9���@�����>[H��_0Vձ!�`�(i3!�`�(i3�&8�,�-��A������t���hQ�GvE#�n�%G2_�ĉ�j!�`�(i3!�`�(i3-��`�p��'v��a\Y������6%�a��<H��c����L�{!�`�(i3!�`�(i3�X;p`�ct�:��RE3z%�u�܆����>[HNl����!�`�(i3!�`�(i3�&8�,��w�Iſ�Κes��O7p�J��PWV����ft���}�k!�`�(i3!�`�(i3�����_��R�)d
ӳk��,�:�N�*�x�s�٩���M�zp�p+!�`�(i3!�`�(i3-��A�1���q�\4L$ֵ�)�ak�m6!�`�(i3!�`�(i3�&8�,�\������������%�����!�`�(i3!�`�(i3!�`�(i34�0 L?�p���@Z"]�ϓM��!�`�(i3!�`�(i3!�`�(i3�X;p`�(������6�5�p��-sx=!�`�(i3!�`�(i3-�����D)������DV(�|�\m�� H%!�!�`�(i3!�`�(i3�&8�,�,�2��E�7�k=��#pa�ǂ�?����-!�`�(i3!�`�(i3!�`�(i3K�1G{K/�t�{#	�x�u��߹c��!�`�(i3!�`�(i3!�`�(i3��%ў׫>V��2G����G!�`�(i3!�`�(i3!�`�(i3�X;p`��_�4�����,�n�en��4;�. �e�v��ҵlo�]�S�*�C�3�%@ra��^Rǅ�L,���eߦ��U�9H\e1E�����(�'���:?���