��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}�����`h�ag����pH��q$.:&R�nU���T��ײ2��>���^k�/7�?1�(�c��ߘ�]��|�G��f�:��#tC��o�Rb�v �mD�?�D��L���_�L�Ȳ�V�溜��D�,�H�9� I�����5O|��N�w	*D���y&�f��+K��[y��ڂb�nP	�'~�e�r:���/lt�3� P�;��1�-���/�_m��37tw�n�&/uP!ߌ��˼�{�&�z(ݲm@�)yH�I@'�ew2�\�蝆�u����l�|���j���BR�[_ň��h��Ev�i<l�e;��+�q=w��;�L���om�Q*���T�K/ZT�@a���V������������d�kⲬ��;�Ӏ���b�
߬J�8`�J{D�9h�@dw.+��CLP� #V���i/������?6z���U�6�����w�������
�8��X
#%QG}��>�����<W,�O��x5w�@mG������aV���&V�J8:I���E��ޙX��}�"���(�TT�c�N���h#�K7���=#�hZ]�*�xŻA7�2 �Q[1I�����w'�\�Q�3M���e�t��yn�	� �x�m��n~�q({L�51��;����'��%Ճ�86���H�aF��6��I���j�r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�E�s��bc�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�yߪm����Y�{'%ssA'����{b�2"��-h|,���(����>S��ә�����/�4�}n'���a*�x���� ��V�h�����^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[n�+�Uz�QL�W*g;X����ˉ�1�:�Ω�s8�R�	�}�����`h�ag����pH��q����h��,��B	hI�ˋ����RUq���@���k��!�`�(i3l0��F��j�2tCH�f����@N�c�B����7!ˏW���:�]�^��'n�^0oa�]��n�=k>K�����D�5�KMӕ�r�����ˇ�[$@�������Wu�m���l�]�s%p�:��d��?��s 3�:��)�[���6!�`�(i3=]A��O�T=�4e=��-������yMK�o�Y�Q�;�Q+�[Z��!�`�(i3���D	��U�l>o��|��س&<��3稿N�g����u�UC٤Y��
�iC!�`�(i3"�,�>E����-��%Mό���.�p�8��7��8�u?��I!�`�(i3c��Et�p�VU��Jp��T�����|��p�G	kp^y!�`�(i3c��Et��q���U��X�=)�H�7M���!�`�(i3��|g�Y�'���Xw�P���w�8Tʈ�Ym�ݡ��1��v�ј�"��Z鎬�������(���]�����|#9����o�t���⍽а"�,�>E����-��%Mό���.Ӂ��̰�!�Xy|�W!�`�(i3c��Et��q���U� бb*	��|	�WI!�`�(i3��|g�Y�'���Xw�������36��T�%G�D��#�]2�y�Z鎬�����	�7 �#֯���, e���TYl���#�]�!����M[��Ǣo;�Ul�|�Ƀ�?PA?e�J$b6�I��w��,c�A�L'#���h����`y���[��N��>&S�XQ� ":��v<�����
L'���Xw��ˣ�X| ���j!�`�(i3�]2�y�Z鎬����(��eظ��6�\�f�!�`�(i3N�By3��<�]�!��	Ǹ�y85���~iI�D;�¬pX��g��U-�e�,���6+��L�t��n!�`�(i3�"B��$I��w��,c�A�L'�iR,��5�%]���a(􆿳����^�����Wj4��⍽а�����E��@IE�U��*�QN����n/�Ǭ�#v0V�b��F�6ѫ-����#uw�Y��k��ı��*���q{?d']la�b��Wa�b����y�E�nwE��S��q�P ڨ���"kA��8Z�ZVq+��T���jB�Fg�Y씤`��p��>�B��7���
�-C:��������*�+w�7�G�6�!~�!�`�(i3�n`5�fK��@5���<ZJ�hEc�>�T��u��!�`�(i3�E����FZ鎬������_�,����XmIOO����&{�Iћ<���d�٣���N N�S�+w�7�7,R��(�ٰ�Ř�hw��z䮃\w��0]b!��u��K�&�a�PB����A���+�J���q���U��@����gG���������g��E����FZ鎬������_�,�;�7���c�5��(�V�5e}�mhU�d�٣���N N�S�qg2�K?\���=ZXR΅;&�_��n`5�fK�\w��0]b!��u� [ad���e���b����+�J���q���U�\P S��;
�i(���ε}R�4�̛����)�~V�G"~��.s��I���:f��9��7h��Fu���!�`�(i3,ԯ���gn0|�>�ɏ��t%>^����80�i�F|��9��a��zr,/�؊�"�D�S�豗a�.�Ӂv�u�o�\�����s�^΁�a�n����I8I����T@a\P S��;
�i(�����ȗ*Zx�eY@�)5�(���{�eV��� dQw��E����F���h���eY@�)5�(���{�eV���C�T��,8�mԘL�kѶ���� �%���ߤ�>��7�4�f�z/1���"�e��Ef&W�]��X>�i�
am�B�홛���=����b��|2�5����`KiW��
�!��E!#�1����8�TP�M��=�&&ĕ^$&��Z|�W3���U���P4ǲ ��� #J�Xh�hk�Ln��S�W�͉�V��-d&�.�_���y�wN���@��}�
�?�$ϙRl�b����aYM��d�٣���N N�S��E �����VF�˷�зq8�Ј'���Xw���,DFmғO�4}v�7b��n`5�fK�\w��0]b!��u��B�+2��O1�Et�]�!����w�Հ��a�e56<�5{ΖM+����+�J���q���U��@����gG����s��p0���Y$�7s�9���o>��l%i�-He�-�c��3E M0�A����2Z鎬������_�,��i�p��+�/s�1��p��Q]� _�rs�i���`�M�	=̞��>��vbëdP��J��@�T�\ ��i3�|)sՀ�i�p��+�P(�s2�Q0���~*��ό���.���K�Q~��\������T��7s�9���o>��l%i�-�ȓ�iӚ/��E/��FH=Y��@����;q�D%���>���U�����:(�� /�o8��N���&U2Q�4:b���n!�uo��8�����JC�� W{�R�$�V�<�`A��_i<tb�N^��MQ���0�E�`JcU����;q��\���S)��y��숕iK�D�b=W�<ish�Ž�Լ^=Г�m�����g��|�;�Ojz���)e��ߧ.�go��1�dQ�����*��� PB����AP�p^� ��X,_�1_����2�K��n@�Xy|�WA�$�����jd�	�!�`�(i3!�`�(i3��+p��qR�D����/uK��zk���Ҷ����S�q��F��L4ߧ��A"�7qz+�XЙMǿI?�3�MO@"��<=
pαL�*
 �%w�*�7��O�Vp��ZD��u���m���d�A�$�����jd�	�!�`�(i3!�`�(i3.��J���8�y)j+| ���j��X�z��p�:��H�f�J��
�fڨ�y4k���Z!�k���Ua�t��]�'3�e�g��ЙMǿI?��d��{x��O>�7�,��n6�o8:4�I���c�90Mj�dL�N}�m��{x��r/�%���$����]�!��	Ǹ�y85�A�'5�i������4��k�y'��a~WGS��yB*��/qRr��G��2�
:���&X(O���I�{u�ݚ��O�������q%��ԏ�:Fa�7����os�鮊��h��<���"sS<GYqcHTX�';��#jhDJ��3ish�Ž�� 4ȶ>~!vk���������|e"��\���S)��p�:��I����~u/��kOT��f�,�k]�<<��%�"�,�>E��dN�<@Iv��nt=:��:5A��p�(R\֎u�D��u�(na��[%��/��kOT��f�,�k]�(�[�*J�a$�Y )P<�ܓ�Yݑ���&�d���%O�	^���y�įէ3!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^%w�*�7��.��Ã���¢	�B�d�ish�Ž�Լ^=Г�m�W���b�0�J���hB;PB����A����;q��\���S)أY_����f�,�k]�<<��%�"�,�>E��6M�Z�i����fd}^��5p�T�ۛ����˨g��U-�ew{�I��!����a�}��l�^!ЙMǿI?RR6��-z��	h��4������l�e>%������)�δ��Iћ<���I����~u=7�7K�PO`�� \)�(R\֎u�J�g�*�)ʁ�]VaaV�h�iA�qIp��K�������;�P�t�5��f�,�k]�[��c�"�e��2�Hb6M�Z�i����fd}^��5p�T�۞�iL�~��\E�W��4b�^�#�n���<��j�z��8��#��)��.���q9+t�}c�n��`Z5Z��k\6�c�
ox7dh�?����k��㕏~�C	����dܟz^���G��B�+2� ���US�������q���f�e�x��w����PB����AP�p^�8!�|!��[렾������z�կg�R�<<�U��x����2�K��n@�Xy|�WA�$����Ҍ5`��T ��(՛Ny�����ȤЭ���V��o5]�Q;�im��ȍry��	b��
ߎ� n2ϒ�ȡ�&Y��V��G8T�w�nf�?ǉ�=��w]��&�4>��K�&Z0Q���s��5�q	�Ɏ�#���?���,�v�q0�~��̚Y�M����4Wt#��wo�V*T�|#HK�����\��w��;�����m�Tƻ¿DĢ�WZ���6%�a�;�.A�ى1�#��d_!�`�(i3�a\;V@|ऩ�jU/�\���WO+�jqh&Σ�h��I�
C���m�o��vPD��<!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3E3����.��FO�&�X�0���X�q!�`�(i3XO����0J�y��*?(�k�+9=@�#=���ix���!�`�(i3��ԫrI�C�i�4��v��$�V��bst�N���!�`�(i3�#ŪS�������k+�r������z�r{]i!�`�(i3�X;p`�*����V3�3z%�u�܆(��.�����R�!�`�(i3r� ��i�(���B��������23Fdr5"�?X}Ax���x��~iM5/�S3 <-���w�E�V{��a�}�$Ϩ�;?���*/�|�-���w�E�V{�?�k�V�?egE�@��i!�`�(i3-��k�I���ިg� a){��Rk��?��q�M�4�a8&N C^�R�)d
ӳk��,�:�N�*�xX�ϣޓ�!�`�(i3�˺�Q�����C�%�Ko��1C$mQ��!�`�(i3B��亁���&�%��Y��j3����(�a��H��bf�?ǉ�=���ٜ�]�X;p`���){��z��l$c��!�`�(i3x�6_s/�)`� ��q/�"����!�G���-��/ӳx���{L,8gf�mk�7�N�-��#l'U:�g[q�vG+|�<A��4�h��T�?Z��$�~c/`L����D:f�?ǉ�=���_͏��X;p`�����G9L�bW�mT(]a%ڔ�&8�,�eVRN&{�GC�蛝p�Ɏ�#���?�5q{! lczZ����P(�s2�Q0�L@]HS�GB�5��&8�,���;p0�Bx�^��n���g9������@������X7