��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�=A���>�L'jf-�6U�P�H�q}��������]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R����h�K�5���� ��1�:�Ω�=A���>�L'jf-�6U�P�H�q}��������]��;�I�����)O��Ξ4�"�\�� ���K�O�{����a�s�O�ET?�(�c\֣�I��B���t��|U|�/֚�?d��Y�Y0V�MG��U�;�\����vg������W�aeYgA���z�Ś��
��H,7f�t�뾌��lr�)OI3��(�!����Y�f��a�Z��V���a�\�nq�M�4�Tڢ�]�
4��`DA�rS>-�O��<$e|����w'��1�:�Ω�=A���>�L'jf-�6U�P�H�q}��������]��;�I�Qg�@zh�S҆�|n��1���Nޤ�YB������h}���U�)���,N��ma)�B��|���{������(��^9?�\�N�u��.tƶ�.,NYD@s�i��) ��c#�k�8���҆�|n����:Vx�p*��� 86!�{��&`;gf�+���h΀��q������>�r�O��C��0���M�<lbts
�m�;�t��q׼'ېoB;sѱE��q�eX;^h���l�a��6��քL�02�|4��?�-W���raУ�����	x]�<��O~����@N?�q)}J�5[�u8t��>䙙J�S7^�	����5�Y�w��:�F'n�//ChR�,��}�Hy�Nk�m����*��O�t;kV�XD&w��0���q�M�4S2��#�;�!_��(0���r� ʢ�p\ט~ٰ�Ř�h^�������;�g���\ۨ���� ��j!�
�:f �k�8���҆�|n������}�K1!�U��ci��j�|}��f�+����4���_Xsp#HXD�5@��=�Ä���
�V[�g��uh������[�_y����]����F��%�����Z��\bI;1:��8&ͽ�m�!=�y����h�}�_nR�� ���E0��^��w�qN��U�)�h���_�[e�t���/ٍoE���dʡ��G�YT~���$mZ��^���/��ʍ]�}��{�ڌ�2�E�= c�J��������+�UZ��T��B���6���k�8���҆�|n���(^k{3�ne�T.jic#��-m�Bf�+���3�_4�j��)I��U����3:�K��9���- J�����59�0O~��P��_ovt��@�m�w�]ݞ��+Q�?f&��7}Wo�ֿ#��L�����RL�a)3���ʉ�Z�o/5�5�R���O����r'KZlֹY���8���+��"B%.�:�*J��¥��1rcܛ� -n��\�4�s��{��]Q��(�Y���m�����h���i}3�L����´�^� �Sr�O��C��0��$�>��w�����N%
��̥㡡�u���;�Թ!o�o,%H�%�p��� ~�/��_� H�C�I-�#��h`���r�O��C��0����bm���?������@�����c�J���<�"F�6x�_uS�CO�����U���o)��W�a������qθx���]8d�\�:H3?��n���N<�n�]��xw��猅
�V[α)j�o�R���V�8yd����Eg�~p!ۓN<E�����@���ަ��%�|%��]
�V[�圉��`�q�r¢w`�&qQ��00�c%���]>�x!����<u��w)�S���f��^@�~篟|�<8�F�-:��ԧN��78�:r&@��$�9��_,n׎ ��73��>g�����Mp᫼���hvK+�va��2鍔�	g\A.����S����9��m�!=�y����h�}Qd�Аrq��;nQ����>o?�M��;]/d^Bg�t��P	�x�[U���zy��<�hV�q��KPi8�����m��d�7������N\Q
7��0���Z�I��y�BR�J��?1;m�!=�y����h�}y(;⟝*#>*��4D�V��(v;o?�M��;]��,��K!�ۻ2�e�1�ΟÈ�bHO���1���RL�a)�Vu~c!�D�-�W�1�H�A�;�q�u���;��I�6r���TJ�2Y�d�To��JCq��jr#�9l$\c!�/`C����G���ϟR��H�<g��ũ��^��Bc��P���3�3Y��P4y JŇ�E4�I�E�-�rd+��Er#�9l$�^����ݧ	�Y�����\�4�s��u�@�
�ԟ�d��c��u!^�8�Co?�M��;]�NT[a��<_��e�ް���
*-=�a�g'�_��z��c�.[K��mN,����0j Oag�1ݷ�NC.��6L����kE�/אo£A0��/�����R��N��:ju��ƴ����RL�a)�ƞ��U<��I�m�$�Z!�e��|�٩7C��H�pc;}ita�Sc&R6�}�t���RL�a)r��fI�����,�%���)0!�Xl��vrǍ���u���;�z-�~	2�O������|�OA�
܊��?Y2���3m�!=�y����h�}jh�6g��+��� ���k�o?�M��;]�Qs`k�sǈY���K��j�r��!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc(#`��Gcp��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�//?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_E$ô&y��ѬL�1m��+Y#_WӇ�s8[ZΑ� �}E+�E$ô&y�y��ά
d9�[l�&��q�©���H��JnXe�+�Uz�QL�W*g;X��'p�@�I�?g�f�ja1�n�[�ެT�Z¤��I^��?�;��XC�_42K�,\ަ�It�k\,آ(&l������g����=l0��F��jT�����N��2�F�PǙ#Y\��?�l~�Uf���}��\�v�T?�7G|`�UxHj,��|��	�"�,�>E����\�v�X�zgq����2��̪U��֜��3"�,�>E����\�vņ�Q�]�ޔiyV�[R�^Ƒ��!�`�(i3JHn��z�_c)���8���bg�1�Z���=�������b9����,����d���z���ߘ�)�I��<
DN�l0��F��j�q	k���A���������]c���H������i�=]A��O�T=�4e=��-f[� ��³��w�[��C��!�`�(i3���D	��U�l>o��|�,+$\�M���j��"n+0�l�R<�q��f�}��Gظ0����!�`�(i3��|g�Y�'���Xw�f�VHF��Q�#<4^��E����F��j��\w��0]�\�LtF�!�`�(i3N�By3��<�]�!����M[��Ǣ�<��>��%@��4��c��Et�Y�{'%s�[�&B�踫g(�r� k�|6�8�3 �;]�F˯�+)�"j���b7|#9����nސ��3���w�@V�"�����/�]�!��M8���	D%��_�ͅ��/��=��K�q�?l�_��Vx�%L��W��_�ړ8���/����R�Jm���S�����*���j�Ƿ�:h�(n�_cn��\N�2߄�2W���R0L�>��0�]2�y�Z鎬�������(���_U)�<�&#R�^Ƒ����"X��[s�o0�` s�"��=�6��w������
L'���Xw s4S�'�i��`�z6/������,���eFz����zf�U����z~��6��	�\�HP@�a%=dϖ�i�@O�x�7���q�©��'w��
�fʖG�œ����s��3�m��L��]�>-iu�`���`�+N��?���&���#�{�0;�}����\Ҥ�Yk"1/р�{:��'��팣+����F�N~Y�9���$1m���0@ȹWpH7���
I@1���t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s��.|Z���I7��-5��6��	���`y�����g�,P�n�Ͱ��Le�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cUL3�X�j�>&�&i�"j���b7|#9�����ѩ<D�n:3M �[e�~'��Vh���*ܑe�W����n�4�{lGD�V�B��иܖ��A�.u�r���,DTc�~y��i�i��욕�'�e��`�)�	�%{�;����f�kN�ı&l����[}�@��L�(��$tI��'��d�uY��dzw⭏l�u��s$y�<5������U��֜��3��P=@��������$��Xo�-��8�%���ތ�1��\�v�?M-��6(uU����z~
������'=����V�Տ���i����_]���T��\�vś��Z1`�<ͯ�G��R'),��`�*@6��8���M���de{���W���g�,P�n�BL�Jx��������k�V�6IWJE�$��dg0J/��=��K�E��{#6�aw�"�HߢI|{�0Lʡ;�¬pX��g��U-�ez�r�6��DP֞ �����Ə�_���ބ6WpH7���
I@1�ؠ&���Z02��`�z��GZ>.�0�i�ܰAb!��u�mj�B��V�}0�z��[��Q�՝�i�(�S��]Q�I����踫g(�r� k�|6�8-+��B�G�
�CӞD��]�)g��E����F�BL�Jx���`t�A~�9�{u�:�髊}���ۋ.�?��u�htGW�PA�;�֋`N&l�����*����s��'>s�a�x��{�6�e���ӯIJ ��`y�����g�,P�n����|!���^��\i�@^7&ģM��i;'~��% &gp�	8���R}�
�?��9�|���l�d�EW_�Բ������5�N�~u�푧)���x��ͯdoP��a�I�;�Մl Q5b11��m����ɨ���0�]cJȷW+`�x�ogJ��S0����~���N/��=��K�����\l�'$9�F<�'a��T���k��$a(􆿳���Qs����� Ei�lmZ,��*�B��	e�2%e"���Z��#6r����I����"�[/�cWM���6����]�]�!����w�Հ�k-p���� <�����;8σq4���s��TaR�^Ƒ����"X��[�z�C���5��_.
ļ��~po硇��;]p^kAO��t�+���LQ���"X��[��Q[R�7}ϼ 8����{pxʟwf�X����cτ����T�=�����ϲ�CyW�f�tR�wX��}�
�?���8�8��/��N���a�x��d�uY�ا�W��_�ړ8���/�a'�<� \�� |+vܽ����#�� �d�٣��c�A�L'�ٙŧ�)#nJ�|m��g��U-�e5��e6²��_�Ps�T��������a��7s�9���o��S8�u�?�f�R���k��$(�%�8���Qs����� Ei�lmZ��x����7A��(�n��rs�i��<�M�AϦ6��.��L�L;Л�����Øf�.�Ӂv��9K±�sR�{F���d�C�R��C�<x�P�$t�[�z9�[�s+�¤]�o"�s�8ĩ�XZ�#J�~5#c��HՋ���)~a���@=������yM����?XW�~a���@=������yM�U���!=UgR� �ұ7���?�!�p��b���A ��2������������(į$?�d���&�/��#X�>�혅vº�w�⽒�k��q��־�W+��W�f� 4�qK��v��z�NFX�5�B�ʏ��Z��PlJ�M�=�혅vº�w�⽒���M��ҹf�f3';��|B���r����R(ǜ`���IX0F�MV�ҁGG�.Mm-;�!�`�(i3��èV!�`�(i3�'ž1�|�'����u��r��!�`�(i3�<��>��h�EtC�<�b_X�XV�b�z'hۉ)��d�7�q�!�`�(i3W����GS�*;q��=<�6>e��0�U+�qbp@�!�`�(i3`���*1
�:qEptiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3�s�Yls��8��GM��-����!�`�(i3q�\E��0�����?uA|�d��?KYC'v�}M�9s��!�`�(i3��.J7h��r��H҆�.A`��x������D�f�6l�}��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3��ܐ�}ħ@�BY����;b�-�2�V��	��y>�����HN��R��?�d���&��g�]Wt~��^�V!��� JO��"�5��Dz�͒�p��e"5�O�%E#Pq�\E��0�����?Fe��1������Ə��}Dq�f�mj�B��V�-vR�Ψ������S,��!�.�g3ZE��g�Hb���KF<�w�R���y�sL]~ц����kUiPO��sY�Y8��t�9G�#,��gR� �ұ+s�Di�R{ZL��틧�gR� �ұ+s�Di�R{LdR�?�9�e�D�a~�'�� 7��
�+�0��H�/zP5�O�%E#P���E?��>ݣK�6<o�����w�_--���gt��,ۛ?ꢰ5��܊S�*;q܋�DKY��,Bp��S���Qѳ$G�;��|B�6�'Z��OG�6<��.ʀ8�t�|2;$�JأͽgF"?�Q��ǺΕ�f�f3'_��s�֙����N/Z�S�޽_�c�{I��L�1p/-�������?�/5��"}�a�x�mj�B��Vh�EtC�<�YT�oT*p��p��&�[���t�T��?E-h��$^(?��"�$y���Td�HzG<<�6�Q=�r$ɓǃl[�Ƶ�1tSjv��� л�=��,���H��nF���<�W�.�P�	��
�Q�}�^{T~H��璓�c�������t �[l;[�G���KlG%��`��ǚ��ظ
��@�U#<�6�Q=y�}�6f&rG��Hb�T�R��!�`�(i3��#
<�(z.Ю;�Ƴ0��atN�s��S�+�ϧ>(Z*��b!�`�(i3��4-劽51�X�c�rs�i��]S���D�'�)�Բc>ݣK�6<o�)�/����O��]��MԵ�x3���ʗ�%oc�����k��u���Ra])n#6�E܂%d	!�`�(i3�/�cLbŪ�����:Y�{'%s��$��S���b�Bϱ��<��>��h�EtC�<�+������L�*dgN;�r��H�?X���V4&�zʖ>��;!�`�(i3��Ě�����}Dq�f�����^���Ú�'nB�Qטg�u2Y��Pv����ʗ�%���6�7gE�s@�@�/�M��C�x���ݚ�Н�烉s)�v�bP�63Z�t��Qѳ$G��A0ok��烉s)�v��IX0F�M0���w�����,�ǰ���!�Ab#��Y��F;�Ř�T09�����\��+x⣗�C���c�)��|ԛ�iP��!Ʃ��J�8����+N��V�/�Eԣ5��)=V�S
����fk�|2;$�JأͽgF"?�Q��ǺΕ�V�܄WD��|�����:�EB�Z5�O�%E#P{y����M�V<�'��zX�k뮏��y�g�e`�!��:U]r\^ؓ������b�� �_&l����}@4���5�O�%E#PZt%��m&<XdYʼل���OH��c���鿋�E~��k}����/C.�L:,�s L�Zl�W��{��]�L���/=9'�����mC.�L:,��i���A��ݚ�Н��9�|���l8�48�{..�Ss�g��+˘\5���jmY�VS���g�n�{�6�e
��>�i�g��+˘\5���jmY��X"e_�4�{�6�em�;���HN��R��?�d���&��Ebu��SENan&�\�0Iѓ�1M� Ѯ&U��8�>r&��U������yf��>5�O�%E#PZt%��m&<XdYʼل���OH��c���鿋�E~��k}����/C.�L:,�s L�Zl�W��{��]�L���/=9'�����mC.�L:,��i���A��ݚ�Н��9�|���l8�48�{..�Ss�g��+˘\5���jmY�VS���g�n�{�6�e
��>�i�g��+˘\5;WT-�bԬ= ��2��' ���@�$� %7䨉��%>�rG6j�"Hs#<�&Ʌ��@��v{�G���ށ��YxƜ��3��O	�T/ k�|6�8�a"�/A$���Z��!�`�(i3��`!�r7��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ����$�����E~��k}����/��&%�:z�+���LQ��:5A��p!q��V���'�Pp̢����{_8�Y��=�}�Vݨ��}Dq�f�����,�ǰE��C$��C�Y�\�P�p��jN˭�ޱB0w����u���ei�j���s��d���!i��'T���+���J�N�#(�����+�F�$-��,'�*;���#�b�PSK=�>���@]��}Dq�f�����o�a�NO�*b ���?R �K7͍��|��W&":�;b�-�2�V��	��y���SM���G=X��t,�K4a���ݣO0��Z6�o8:4�I���c�90�Ǘa��xO.C��|#HK��A(�c���_G��Hb� h�ҩ�!q��V���$��v�ag��Se��0�U+�qbp@�.�x�BEVݲXHBB;�T�dN�<@Iv��nt=:��:5A��p��$���͜P_�_S:g�RMm�o��'����N��U��;y��v��\���
^�ݚ�Н�y�}�6f&rG��Hb� h�ҩ�SƏw0���iD.l^S�ñ��̞�9�|���l8�48�{.z�X
3kZ���8�q����1�t(U�l�XdYʼل��OY'���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�Mt,�K4a���({�Z�f�q���ۈ��J�a��?�d���&�ϪE�smy~�K���@�{�f%���s��e�i��B0��J����M�!�y:i����2�x�h������M�!��^��BcƍItJm�Ԗ�Б�����ph�)�s\Hn��;��|B���r������/��r3���ҕqC�G����]'\gWg��	�Z�kfc&�2����ʃK�,��`U��B��-%G��^���j�VD"������� л��'ž1�|�'����u��r��<�6�Q=��hY-N�g(�����x����E2b�z'hۉ)��d�7�q�!�`�(i3�ٻY84����<	s/����AIe��0�U+�qbp@�!�`�(i3��b��~�F�KD�Vr[/}>5��0�B� �b��!�`�(i3��fCI��8��GM��-����!�`�(i3R���Xc�Q�R���F�(|��8����ei�B� �b��!�`�(i3�� л�U�~�vmȋ���OH��c���鿋�E~��k}����/C.�L:,�s L�Zl�W��{��]�L���/=9'�����mC.�L:,��i���A��ݚ�Н����y��lDU�n�X��zq����1S�Д_9[�l��a+Ĳ
�),��Tt�j� �"�m���rwӷ9J�E[�l��a+Ĳ
�),�5C��-��"�m���r!|�α+!�`�(i3,�u�S�v��T/q3b�5*s6=��GZ>.�0'j�j�Jy1tSjv�!�`�(i3�B�.�4Ӭ�P8��PS~�Dn��i�Q׭n�L���/=9j���)��Q��\@
��:�)�<�����⪂!t-�u	D�&���A3�Q��\@
����G3҇
!�`�(i3�� л�U�~�vmȋ��OY'���c���鿋�E~��k}����/]P�����+���LQ��:5A��p���y��lD�`6X��gO .��0w����u���ei�@�ܫ՞�� h�ҩ�!�`�(i3�iڈ(��֟�z��n�*�&�v������⪂!t-�u	D�&��9o�d�E�"�m���rwӷ9J�E[�l��a+Ĳ
�),�#�T��6�"�m���r!|�α+!�`�(i3�B�.�4Ӭ�P8��PS~B;�T�dN�<@Iv��nt=:��:5A��p���y��lD�A�s�d�!�`�(i3�� л�U�~�vmȋ���OH��c���鿋�E~��k}����/C.�L:,��i���A��ݚ�Н����y��lDU�n�X��zq����1>� {�}���my$�N��o�/���;!�`�(i30��l!���O�D mWN!�`�(i3��&.��8�F�S�1 �0��l!���O�D mWN��\ Nh$�)�vx%�уZw3���ҕqR�<�t@R��X鷴QW�w��fD^����+���F�}қ~�C탤ϻ�U��)���Y;e�iKI/B޾PԐ#��go`iI9�o��|#HK��A(�c���_G��Hb� h�ҩ�!q��V��hiLi?b_X�XV�b�z'hۉ)��d�7�qĹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv���H�����Yu�������&G!�`�(i3�9�|���l�T�3#��6��:[+b��$��v�@���BEVݲXHB��Q���N�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��jr��*�t�1P��s^���dm��\4��|�]�+M�6��cb�z˪�y��?�w-�G� I���~=����M����V�܄WD��|���85HF���h����,�RVo)MP/���:��9eɽF�	?�Ľ�`���ʰ�c��D�C���,���Ъ���\�rҖ�A$�P������5d�`UNP�{y����:�*" �`�r$ɓǃl[�Ƶ�1tSjv�SƏw0��,��*�B�JQ�jƂ�nF���<�W�.�P�	��
�Q�}�k��^�1Aj��t�35L��$
8��2�ֈe�cN�0��ž�Ć�T���7X���c�}��
�t��T&���LQ�/81tSjv���'T���+Ho}2b<��8�.-M֑�3����H:H;��G�� O^_'&�d�'fU����"��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M�"v�(=�@� �-k��!�ˢ6j�"Hs��'���5W��1ReC����&rgG�I�4~��J�O�R�[P�3Q)ъo�Ʊ�_�eD�Iѭ���N���c7�t�~�<ͯ�G��R'),��`�ӑs�<`����Ƶ��U��R�~z��	(�L�������Ʊ�_�eD�Iѣὗ�L���#g�k���:��Ɂ�]�'߭`��@_��M���o��_�Rv�䩲$���dS@Ɵ�od�G}%��b�l)�=����"sS<�0�zG�������&G��'T���+Ho}2b<��8�.-Mb_X�XV�b�z'hۉ)��d�7�qĹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv���H�����Yu�������&G!�`�(i3���JQ����c�0�=�8�tw��~~!"s�x:�^{ʓ��ṵ�0�)!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��jr��*�tZ�u�x�c���2c�aI�FǤF5U�?�d���&��֟������cI�M�A�E ޴�g��.���f��Pޤ��I�l<�*X�M�m��B&�� �=�3ǎ��������φ��~�����G�٘��������a�o�ax4]Y����iZ6�w����k�k�V���ֶB�M�K~�L
��?��C�K`bX)>��v�k��}^ZM%FW^AΉ�aխ*>�Ƣ��}K�����ncj��#x������.��4�F1���l혡˘�k���)�Տ���i��}��g�'[�O����� ����H�ʱˡ�^���?�d���&�̬���	p��D�(L�IԬ6`��V�������Hf2�Г�P)��|�"�/�0�T���}��&%�c�J�%�Kw	�FD@s�i��/lns���>}�����L��Ay46�o8:4�I���c�90�Ǘa��xO.C��WHe�Q\���F�`yx�>�+X�M?��y�!�`�(i3_'&�d�'f�S�bH�@>�ö,�K7͍��|��W&":r(�z\���M������)��nF���<�W�.�P�	��
�Q�}�k��^�1Aj��t�35L��$
8��2�ֈe�cN�0��ž�Ć�T���7X���c�}��
�t��T&���LQ�/81tSjv���'T���+Ho}2b<�TC��G�KI�R�''���Xw�j�7��_'&�d�'fU����"��9x��p�5��/��8���/�z�X
3kZ��ɮ������~��:�Y�{'%s	Hu�L	�~~!"s���X����k6��.��L�=��gr(Ƭ�:<��j!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��jr��*�tZ�u�x�c���2c�aI	�U˾���\�Q��4b&��K����G�_���J���Z&��i1�F�\��ۧ孡4���H�W�_�x�l��1:�N�*�xX�����p��X�6��.��L���犑e�A�T�g�v�����.o�%L(\Ӧ�ݡs��������B��1Ʌ�Mi��팣+��9&��)�ꢤ�OgE����T���ɮ����A�����J� ���]����b=���9��稕�a�/!O��8�i(n�
e�3+{�i�m�T��q�\E��0����9!{����*�;�C�kP��>A	�U˾����팣+���Q��ǺΕ�V�܄WD��|�����l��	�?n�@���x�����I��>��V��	��y���"��l�*>�Ƣ��}K�j����wV�W�Z������;��|B�%����3��!S�v?��*&i-1D��VhT��z�,��6��.��L�L;Л���TR5G�!�OTo�aT��E,��a,�_'&�d�'fi����]��E�g�������(ӈ���\��Z�ܼCI�_���q9+t�}
�0���U!�l.T��=9a�Fc��;��i��5�%]���a(􆿳�cof��7��ܼCI�_��Zz�U��W�� ��! ԝE����E2�>&�&i�"j���b7�TR5G�!�OTo�aT��l�^ �p�Q(1CU�m��e�� &mjR}��Ɲ,]�eT�?�d���&�gb3������?��;!��5ܲ�yM<�����;�	�m�`B��ʍ�ca��˛�;��|Bd�SF�v�%��6<jsrCm�k��jiBy�D�rs�i��r�����^{ʓ����-�����<ͯ�G��R'),��`�}�8��f�FX���v�\�b�U4��\w��˪?�-���ei�^�̷ؠJ��:����}V�)c�`j�Txk^��]��3R��������Vo[���˚����Z���2��}�������Ə�m1�ؓ� ,��rQ3���w�@VeX�P�+$r�t�}iV��	��y�� �P�qN#?
]w<�h��R��e�j�Txk^�a���~6�z�����ϲ��Vo[���˚����Z�ם�.J7h��r��H�v@W��}�������D3���w�@V��B|_��j$r�t�}iV��	��y�� �P�qNy�WE~�YV��	��y�2B��$�yuk7�'��G3#uV��rU�w�⽒��8�>r&��H�ʱˡaf)��;��|Bc^���Hp�T82g��	��#�^�y�j�˗ߘ�)�I�����v�h�g��U-�e a⣃_B7�}�!��T��a⨯�`j3���Fm�b�vA`v@񴱝�P���Q�烉s)�v�?�d���&�p�T82g|��!l뜗��,�ǰ� Ϳ�&�vDv�}˨��'��*���E.t�