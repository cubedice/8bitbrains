��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}�����`h�ag������T�h��~�a.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I��7��_�L_H��Y씤`��p�eh���w1�I�?g�f���\X�<����8��U��Ĭ���^W��C*z�w4G�� ��d�n}K-J��K��z������3�z�ω���D���+�	���lF72��{L�8br�.�/�d�������4�;(�GoAW�~.8%D.��n�P��<���-ZW�k%u�e<��⪘����t�켻�S���c, '�yN�210�|��1�@��cOL`¸[
ϊdl�E���2Ee�Y�R2
�I.��	���
��i�S��/��5[��̔��o�^���~�CxT�Z4Y3>���~�)A�t�ە�.U��B�?���@���%M����@�]"��~Ǣ�)�5�d���u>\!����G��4j���I.B�
m�Id��D��4�Y ����Α(���NZ�A�!�%���?#�+)5Y 3�oGJ�#���S��Bm�4��k`'&Bc &�� �~�c��t-߱�~����|��d��^Ӛ�z�?"	��k�8���҆�|n���f�S�z���hݜ�!Z1��,�'��c�s�F@�4%�s	��4�7�t��q���ʞC�ݢ��j�r�
� �AH���g���	�e��ME
py���jF�ۣ��M���F@�4%�����^)�D���%�d��;�
Ҷ�8�U��]>��D�,�Hr�O��C��0��$�>��w���(bV8m�G.]�7�F�u���;��V\Bh���dM�+���^����8M���:\���n�x`��{Mїa�HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0- ��Ckӏ�^!�|�Ƅe�k��'p�@�I�?g�f���\X�<����8��U��Ĭ���^W��C�9���$1m��w�Z�M�_F�k-�!�`�(i3!�`�(i3c��Et��q���U����?�@�|+l~�8!�`�(i3��|g�Y�'���Xw�����U�ЂDa��(���o�d�!�`�(i3��|g�Y�'���Xw��������P���Qi!�`�(i3v�ј�"��Z鎬�����	�7 �#Z��M��
�	^���yN�By3��<�]�!��	Ǹ�y85�����F�>R�wX���D������^́|�A!�`�(i3c��Et��q���U�[��N�������l�x�f7﹏��|g�Y�'���Xw��+x�r�2�6�d�f!�`�(i3v�ј�"��Z鎬�����X���*�����:(�L��%�U�Yl���#�]�!����M[��Ǣ[��l�,1B��CSk�"B��$I��w��,>����C��(R\֎u�J�g�*o3��Y߁t@IE�U����S8�bM� 2)G��8���/���E�d��",oMG~�Յ$�O&��]2�y�Z鎬�����	�7 �#��i|�l5R!�`�(i3Yl���#�]�!���D��L#���W���ͽ�ʇTf�\kJ���I�?g�f���\X�<����8��U��Ĭ���^W��CQ��ņD^�NË�����8�9Ѽã� Oag��Ц��#�"�Q:�{�1k�ZV"���:��#tC���,?a��Q\�_q-�㰻������*�+w�7�G�6�!~�"�,�>E���]�!����-ዧ�[�����bp���Q0�!�`�(i3�d�٣���N N�S�	�:-!@xNm���d�0x�梧���]�!����w�Հ�(.V��������lz|���~{�Z鎬������_�,��LE-L [_1�f���зq8�Ј'���XwI�&�\�+1���}x*ؐӘ��b����/�:�3�TF
%$�����!���d!�O��1��2�.w[�%�!�`�(i3�i3<�f�D.`�Z���L5ӥ���98�
x�?�����tz|���~{�kѶ���� ۹;EtS<FۈJ��R�Ws�N"T8�zn6�u���Q0�lC��ۺ_~5�Ǫ��I�&�\�+1���}xe�4޸5b+�����50)�}�����T��.��W����"�,�>E��ۦ� ~�p�+�����50)�}�����T��.��W�������E���b!��u�PQ�>\Ճ�I��b-���q�[���QR�hǬ�&Q���5r���$:��8ڇ�ȓ�iӚ/��E/��Fv��a���7��Z�/�Nc�?&3�7-��ԡ6���9�̪=����\���S)��y��숕iK�D�b=?#�ˏk����0��G��e���������6~��2��,u��T�KKnfO����&{���x)�o/�1_����2�K��n@�Xy|�WA�$�����jd�	�!�`�(i3!�`�(i3��+p��qR�Ovc�[��l�,1B��CSk�_�#g� |y��$ŧ���`3���jO����&{���x)�o/�1_���_��.)<��O����&{�6�LbE���jVѭ@!�`�(i3!�`�(i3�%ؙ,{F�2�����w$�Q!9Z;<�O��gC����hj���hɝ(z�ZI~,|,���pq�vأ�U�[�m��U��)���Y;e�iK-pm!9�>��n4s1�U��B��-|k������������r$ɓǉ�.y�U=������&G�7���������U���g�'�^����x��7�֕iK�D�b=��p�:��D9��ɰ���|e"��)�δ��Iћ<���I����~u���NM���(@X~�H:������宦%��s��u"���ܹ߆�p�h��d��JXl'�T��~��Uг�|<����&��m���d��(�[�*0��d`��������x��7�֕iK�D�b=��p�:�S1�ӿ�Q�ЙMǿI?����[jMQ���0���g�����;q	�%��6�W���b�0��%t̓�@�8��"�7ό.R��x��� ��2�w����:��q��5ߧE4��Fr��j�|��۞ͤR*̮؂���@������X7