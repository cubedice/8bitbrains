��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�յ�'�)���Ҷt������5O|�7x��������&�ǝ�+zA��]��~ا@H;�W ��W�5�k�s����F��W��`��q�©���?��P>����M7\F���r��C>C�݂�N$��/���	�0���'v6�o�"c����A�&�8d�v��x�۔7�D��:�b�#�Bn	����I@beB��H��>I��4��u"%�������j)j*[��HMi.��>��'��E����F�A�y]M���y�.!/�1 T�V	�tL��	�<�A�}Q�� �P�_ߠxR�	�$F5��wx0�<����O4��X��m�� N�X1јds£����&��ea�8����'�����$.:&R�nU���T�����\�4�sW c`k��M��RwM���	ɭ8�i�p&�K��~�MUs ��?�L(	���&�Ll�ݍb�e����K��U�d?p�._q�l�2����v�`��H6�[	�V�D��~���pKJ�)6�X�e��D��8wɦU��D��)�.I�z���{����V���	x]́��D�F���S�V��Fč�y"3��
f��:�%�+M��m}os֮7�"P3��_� H�C�I-�#��h`���r�O��C��0��`�R&.1� 0��]��Ֆ6%n8��u���;���A��j`��'�����`U+n%K)��k��Ǣ���N�y�Yc���;��sD���L��+�Uz�QLQM��S�O?�4�ʗ
� �AH�T�t��3��e��ME
^����c�:���0�F@�4%�u�L�r��3�jT!�K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s��e�IC�_�\H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���%	v3����Ms�JFAa��Bzb;ym��+r��JʅqNA��d��1�:�Ω��
�/�r��]���P��`�.�D���J7"���`���lY�y��
r�(����5�����x%~Y�1�:�Ω�S�T�;Ϗk[�^��_E$ô&y�ݜ�&�0�-h|,����-�KJ�訄��ˉ�1�:�Ω�յ�'�)���Ҷt��_42K�,\ަ�It�k\,آ(��XK��(ڷ|��'�u�'n�^0o��~+�ݗ����Kp&�@���k��l0��F��jT�����N��3w:��O%��<������4];ˍH�F�� g���t�&_���9��E����F�'n�^0o��ҕƦn+0�l�R<�q��f�}��?��[�<��z��}�\w��0]Y��
�iC�o��C!T*�q���U�&��GE<�N�By3��<Z鎬����(��eظ��7�
BcyMu򔲊'���Xw s4S�'�i��`�z��4�+|'Tԕ���ߋI7��-5��6��	���`y����ꢤ�Og�?�#B,�Ң�{l�f|�m�jp=�>��o�
�v�ξ����LUG���>��Oޏ��F˯�+)�"j���b7|#9���{k�h�++k&v�Iz7G#+�ǚ'b�t	�U���C��O]r�<Uee�,��3�L���&Ã�M�R�^Ƒ�Өg��U-�eaԗ5��C�6�ǌ�lA�1�:�Ω�յ�'�)���Ҷt�~��`o��0���r��X/��4�q�:�"��yȯS���Qߵs<��7�m��+ r���7�����|c��c!9M�؀qjZ���A3�(N��㎏qló��|�����V��ߝD9�{��灊�O�i���Z鎬�������(���`$�P.eE���lC��U�T�\ ��y�.�`L�/(f�|��*ܑe�W����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�����څ���D���J��8���/�I����"��T:���V�|�%�|>��A3�(N��㎏qló��@d��שt�v��I�`2ڻ�Ϊi3�|)sՀ�T:���V������!/��A3�(N��㎏qló��@d��שt�v��I�`2ڻ�Ϊi3�|)sՀ�T:���V�#���9A7<���������	N^�U{xN��i>r�<Uee�,��3�L��-+��B�G�@����gG��V��#wFE����_|*uN�wHZr��AR1<]Q�I����踫g(�r��!9nV�[}�@��L}�
�?���J��s�D� �o��z*���Be�2l��4��a��se�ξ����LUG����i�ܰAb!��u�
8�<ua�>����׌7<���������	N^�U{xN��i>r�<Uee�,��3�L��P�Ɏ[`b4�6@|�.�xhf�JF=��,��u�Y�KG�ξ����LUG���E�����+T5�O�%E#P"K���BmY?H/�]�!��	Ǹ�y85�K]���j쮃'�)�Բc�92��4��}�<��}�GvȻ9DO/�rs�i�gsf��"ȳ���u(:h�����*x����[��Z��E��3?�d���&�= +i�1���+�T[nq��ތ<|���ZiXQp�3Y#�踫g(�r��!9nV��#W�U��ظ�d���!ia���ž�����U�p�[���������
�N���7�}�!��+�TM`�ON8]�؊���51�X�c�rs�i��]S���D�'�)�Բc٥\:�l����#w�mc1s�B�~����(��5L�*F��!9nV�ܢ���E��٥���E�i�m}66j�"HsEһ��g�.@�y�T�$f`ƴ��4S-(s����Z$�j]x�7c�oW�Rd���=�W+��W����f�Rs}
#����P�D����Y�{'%s��v�9˞�]v1�_ُ<�1sV�[[��}�.���pqo�}�I����&��Oq���4�+|'9�	M������#w�m$r�t�}iV��	��y`�a�W����u/A3ʅ.�g3Z�`�e�%R<��d{ӆ��^�p~z�r,Q17�b�����d���!i�!�Ì��_���މ��~H��bωJ�³5����XK��(��s�Ӻ���?�d���&��;b�-�2�������A$�P������5d�`UNP�d=��¾ȼ!�`�(i3�'ž1�|�'����u��r���2��}��ăz��r��?r$��K7͍��|��W&":�ݚ�Н�*qA����6\�4�@�� �-j�1tSjv�����l��=�O�-v�*_�mS8<�n�ݚ�Н�?V��j�c{����҈#��: x��XC��F~z�&�?:,5�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ��׹��4}4H��}�	76�&�;��|B&g�r,�2'��;_��8W�w��fD���+C�!-��x�� O���ƫg�Tn�\��B\u;��|B6ϔO��)��Y.!�iɼvA�a�(�.�g3ZB�ek�5W1��g�QB*yT���j(&
M�K;��%YM�	�v�3��!9nV܁�8y�Ɋ����Z���F%�X�����#�݁�ƫ�P�A�I7��-55x|���MM
��,=?�d���&�t�{#	�x����л����[XP��p�����ָ$�/�x���2��}��H�\�(�����t��P�3�pVK���ʥ}cG���I��)���W�w��fDV��	0��.�g3ZE��g�Hb麭�H�κ'��G3#uV��rU�w�⽒��8�>r&�,��3�L����:�EB�Z�w��"\He�F%�X��k��o������"O��`$�P.eE��o��1��MM
��,=?�d���&�t�{#	�x�jsrCm�k�:��=#��9f2Pih{Ø�F�HN��R��?�d���&�p�T82g�{�Bͳ��;��|B�1�A���^<��\�<;2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���+�~c(�
���P�����7D㒅��D!�(9�#�_o΃��Ҕ;	ۓ��}xF@����?pj����eG�eB�c�*��Ɣ����&lNj���!����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڇ��L2�j{�'ĨuMŃ�,��)��5�fL��
nЯ�O�!�`�(i3D�c=p�4b8��K��l~�(��j��ݚ�Н������L�	f퀔���἗jc��{��sۍ�s�*��ф|�P�Y�����TKP�ρ��8e��}I`�翹,�)yD�KjqVe�Xlf�"�
;���?q�����]�w9"xy�b�G2�d���,�|�7����c