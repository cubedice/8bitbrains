��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����Q%b<Y�D�L|�w.j��6��H4ي��2_)��:B!�b�ؐ:�{T�{df;���a,�Q��Կj��_�L��o¸���Pq����w�Y��k��ı����~K�%��������/N<��;��� B]�pE���	x]̃Dj#^Da����M�$����o��I�绯�t�z����)�,�˛D��w���旴4w�1����h���������$[L���Fj�Az���JU�e��Q]�z]�����X".��>��'��E����F��#�xn��Ӊ���@ -h��7�A����А��䬣��x�Mi��Zߧl4���0�?�1~�x�c&	��/v�&����?@��(k��yg��$]B�ʇ8[�r��xmܵs�����G�9*3�-�&�Uxۤ�(���.X?��M���^����S���	;�e���̇���S�q� P�*���k� ]�Լ�c�,ҹ�$�I`'2�=���gb[�,�#f"�:Mz��ʚF���Q�������\�g��5�=?�/JͿ�>@Qթ�����Y��NE,���fea�H��pw����㰑j�ȑt�b��M
���&�F�P�(�-w���8�aňhinOL�T�o���&AdN��Y&O�EbƘ/�D����~��_+|�ntzhn5T⢉�y{�U��:�,��+��kyf%���G�ϠE{ �W�B�l𛗲k��˿�(�v�)�̎����T�z�)��2n�yw��G�!���d��mc�{$W��%�7��.�N� �򢠢P[�$-��aJl5澙պY�l��"`&c�'N�j��6=�[�D����\�Y�&[R���b�m�鴡`ė�G�2(ٝzz)Kn�P?�����pB�o��$�m]�fB�f1I�����w'�\�Q�3M���e�t��yn�	� �x�m��n~�q({L�51��;����'��%Ճ�86���H�aF��6��I���j�r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�E�s��bc�Ѽ?��Q2�=W�֯�^��N�&��^˻f��sKJ�l�i��p�7��Z鎬����@�Q�2��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i��I�?g�f{*n/�,傴����'SR����.�}|��ι%9T��7����+�Uz�QL<(�P[H�������'SR����.�}|��ι%9M��j@�����nEAJ_�'��P9~09h�i�k1i�f1?�e�Bw�M�?_W�\I���A#|��[�m���w��L�����'�@���,������0��D��L���_�L����\�Q�������W|�.ҨwɷY_GH�7����]n���E����F�Z�>)��p40�zɈ4X"��D�����ˇ ���3�ҺIÙ=�H*.�PS����vbëdP��]n���b9����r*�^�	�M�8Z�XPt.�!ŀ���g��ȝ�0����k�

gY{�o��eId�U�mu�!�`�(i3!�`�(i3!�`�(i3!�`�(i3O�^`Yk	�o%^�G@�w ��hk.�BY?�%�j���p|�4�f�5/�`g4�,�W%JHn��z���o�K�v��Ug�B�z������4-r��|ڑ�H���o���&�t.�}����F�Q���6zJ�%�撁cFẶ��Ϊ���E`�=PEoY��gνp�~Lܮ�G��C�(!���d˖*�t���Xswj!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=�Ea�7��m�]|Y2���L�3GA�\.�
��ڃ�"��E����F���8�TP����������s	IB�;�5�}�]����E����F���8�TP���{��XT}u��Q��WI~�Ct���?�!�`�(i3Y%T��BPe.��xu	�>��l%i�-��E/��FzM#��m�v�ј�"��Z鎬����A��:6])2�����Vc2�����Vc߶�z7��Zr
�0�M�yObFT+V��퇇М1!�`�(i3�����
L'���Xw�j�7���5�%]���a(􆿳����^��/$�ߺ��]��pZ�ì��|g�Y�'���Xw靤�:��D)Q7����H�N���,�t��0Q!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�wx����ހ��g�R����!���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��
��`�VL�f{����߹�_|뷦R3��\���S)| ���j�����
L'���Xw�7��0�$�E�#s�@ҡ?��'o�}a�C��ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�uk�+ȭY&�;���dV���f����"�!T�J�g�*��/�p,��(�
t��Y�{'%s2�ew�a(􆿳��_�"ۆ�-:���h��g5]��C�
�b�s�P&"��>����!�`�(i3!�`�(i3!�`�(i3!�`�(i3&�sw'%�I���Pq/{����I����H��6Xk�scX{�X!,!�`�(i3!�`�(i3!�`�(i3!�`�(i3n���[ �p�ø��.��Ӡ�)�6��}�R�#��U_�������y�!�`�(i3��(�
t�ژq���U�Y�4Eb����"-�&<1����Y�e6�!s}6,o�}a�C�Ǐ˨�g��!�`�(i3!�`�(i3!�`�(i3!�`�(i3�5#<Z�D���� aV��w<����=��85?��k�*�1!�J�G��`�B7dԘ]2�y�Z鎬����s(Ǳ���:����v����	N.s���� �"���%a<��A��r�I�!�`�(i3!�`�(i3!�`�(i3!�`�(i3W�%kԒ�Peŋ�-�Shc,Ϸ�Kr%u���G>P���t�td���52�����Vc2�����Vcb{�o��Ш�G��g� ��^�5��^	QW�Q!r֯���,���j*(xI��w��,�$u$Yo�K�d�$;��(D��2G��
bH~��`��|��f�!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=[��l�,1B��CSkkѶ���� �TnX�g^	QW�Q!r�ԬQ�������ս��]���>����C�������PB<�L�V_��|g�Y�'���Xw�j�7���5�%]���a(􆿳����^��������P:�rQRт��|g�Y�'���Xw�����C���V9{)���ևAY%T��BPe.��xu	�L$�����//��kOT������PghR�P��|g�Y�'���Xw�j�7��a(􆿳�*Տ�*9hLx��UQ�`
Iܩ@�R���!�`�(i3!�`�(i3!�`�(i3!�`�(i3$w�����=��bv.�]�Ⳇk��8�?)���O��+Y#��6�SԎ6�r ]���f�+��T���jB�Fg�Y씤`��p�܂aQ��
~�d�9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6�D��L���_�L����\�Q�������W|�.Ҩ�B�g��@E�f�,,�2��3!kq=���� ��|x���&R��(Z�,��F��s�eШ,W��Ou57���ڛQվ���>\L����2�P왣�Oއ�?tee$[���m�m�˭;{o��n�(Z�ɽE����S�Y���&Y'�Y��#�ć5����`K�.�����?�^"4/���1#��Z�����XP�����w�K�� �ӗ4 :��	��h1��'�t��5����`KiW��
�!��6t�.�=]A��O�T=�4e=��-tE��gVB�3?��}�ߒ�^���P���:����sC�^�+r��[��eئ�=ߙ�@�1�˓JHn��z���|��Aו{$�3~��E/2L#�A%��@���_����'m�|g�~p!ۓ�����+�@K��Np�m~|��SۅV̶�pG|t�L7�����Z�zL͊�q��)"������6�Yyk��1��Rk��?��q�M�4�����F�J]�j�j�DS�׭ԘI��'��>=�[b.|�^��
�>IÙ=�H��`������a�V�Ih�Ŗ���H�G3�c���V?*��4!Х��m��_=�|����dlmS�6b!��u�g�G��0���V����P�n�lx�k��V�4����,D������à�w�`L�ekOF�T��ZBi�mR!.<ή�$��DP֞ "[�GVg!�`�(i3�d�٣���o��D���/h�5�G�Gt�5�GR\-���
(���Q]� _ό���.��7�b����U�m#j[�ߏ����ζ}̤�Z鎬������_�,�/�n�*������˃�I�E����FZ鎬������_�,�]^U�*�!�*of�����E����FZ鎬������_�,�]^U�*�!�e���b��E����FAԢ�a\蟶:���U��^"4/����k�z�I/���`y����@����gG�m�D4>�#���nU�4��X�uʡBs=�b!��u��K��I/N#~8"�Z��H>+�w�\w��0]b!��uፆJ�g�*����3���n`5�fK��0z�cUL�I��6���T�\ ��i3�|)sՀs�?�6 ^��	^���y
�@R	~��Z鎬�������(���/��A����Q[R�7�_+H�]��^���+| � �Xz��⸲��+�J���q���U��@����gG2^o�!�!H�N(�g���������q���U��@����gG2^o�!�3�{~��u���������q���U��˞�Bx$�Z�0�8�>�}�"�,�>E���]�!���e��Ƥ�����bpvuD畆!�`�(i3�n`5�fK�'�&UoPqqg2�K?\z��l��6�'n�^0o**�ХM
�?��j�$����ˇ��t| ��aݓ��E�v���bQ</���/�u7s�9���o>��l%i�-He�-�c��R:k�ڛ)�{� �"7s�9���o>��l%i�-He�-�c��R:k�ڛ���X|x���Q]� _ό���.��7�b����FmғO�4}pi��M0q�0V�ʦ�A'���Xw���,DFmғO�4}~n���,aзq8�Ј'���Xw�Y�r�7"���a�e56<��3c�.����uhP���]�!���e��ƤHe�-�c^Xp�ђ�!�`�(i37s�9���o>��l%i�-�u��Y'G�sp3�K�K�7���'���Xw���,D��=�!�7y�<.��2-7s�9���o;�ƀ�'͚}�
�?��_�^�]_��S^J�Z�d�٣��4�5_�o0b!��u��΁M�$���������V�]�!��"��C������_zx�˔Y�|�8�n`5�fK�\w��0]b!��u�֒���\����	��ܘq���U��e�GZ���i�p��+�FJ�9��V�E����FZ鎬������_�,��i�p��+˫���[�D�g-C�#��RZ鎬������_�,��i�p��+�/s�1��p���+�J��Y�{'%s�:�f~=g(���B���������a�V�Ih��"u�����$<g��g��U-�e�����$VHe�-�c��3E M0��G��7s�9���o>��l%i�-�_+H�]������}�1�#��d_��Q]� _�rs�i��s�٭���lC��U�T�\ ��i3�|)sՀ� ʔ.te`�!���;:=ȟ�H�Z鎬�������(���Jם����"X��[��Q[R�7��B�D�F �����=�#����=�7s�9���o>��l%i�-��B�D�F �����=�Ql��u�7s�9���o>��l%i�-5�e`��9S�n�(�a�/��$ʖT7s�9���o>��l%i�-5�e`��9S�n�(�aް�l��7s�9���o>��l%i�-He�-�cI�؉Pj��O" w�7s�9���o��S8��y�)xʔ�1�^q��1��`y����@����gG��d5C[�[_�Qf%u����+�J��Y�{'%s�Ǹ2���$�mo�6L�g��U-�e,%�0g���l������o��0��7"�,�>E���]�!��8�$LQ���	�:-!@xN�/N���nS�dB��Lsk��c��U���q�
����5�e`��9;�������w�`L��Q8r�#�k&�o��E�
���@c
�}�
�?���\���S)�~*a;ɘq���U��@����gG5mv<rdT�'��L���H��̣��7s�9���o>��l%i�-�_+H�]��o�f��ʑ�?��9)7s�9���o>��l%i�-�
�CӞDIi��6Z߯���ߍA���N6n��nL*Y��w���+���$s�>Φꁲ����3f�{t��uC��m���i2J��K����=�#����=��ܮ2�k�'�����Щ��O��+�pʷ���H�2^�/3!�`�(i3!�`�(i3{�d"����f��Vq�m���d�Cw�Hm��p�@OM.Ir㻧���o����A�r��Uj�z]k�M �cJ$���xQ�1���~!�`�(i3!�`�(i3�>d�g�K�R����\R��T;jZ��*��x���aF<��[��CCQ17�b�����d���!i\o�LCd�$zv�+K�ވQ�:��d�٣�����c����յ[+8�������PX6و�cµ��%��(����e_�b�'�wJ::)!�1%�@�	^���y�Cn�BM߯��
N���Ƀ�?PA%�G�Q�W�C�4M/�S�@9m����1�ܮ2�k�w'�2�P�����p���W�,�_sI�^$D���@��( ���M/*�3���K���(�`�2!�`�(i3!�`�(i3��ɑ��G�:I�#��{����h��N�M�0��F{�r��졾�g��[��o}����g�G��0b��K���g��;�!�`�(i3!�`�(i3�>d�g�K�o�t�����%����	���
�ƫIX0F�MH����M�-�F6}����!�qgjQ�f$~�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�K��I/�@t��U���~=�L�����3���G�k�a���!�qg1>O�^�p�`���φ��<�6�U�7˖�ɳ
xM�v.��ѷn＇�5�v��cg̖UB�nojL]�T!R�ʁ���Mյ���ݑ��3��Y$�M`�K)��v�:�-22�v%��v��!�`�(i3,�˳�*C�����p���W�,�_sa��o���H�RtV�^����&��r��졾�g�Y�٩�����ݚ�Н���w�w:�!�`�(i3��Aڬ&W�����=��w)��
=I�^$D���������P�íN=]8k��.ͥ�H�RtV�^!�`�(i3�<@���ل=����h���}�%Dܭ��}Dq�f�՝� s�#��qX7'��֯���,�ۿ���L��:����iW3��OEʨ�`N/������&G!�`�(i3�7����������EN.74/������.ݍ|�!�`�(i3�̢k���������P�꠼*d�m�d��-��!duP���2
�M����d9=���u��r��!�`�(i3h5���=�t���_j���Gƻ��������[j!�`�(i3��\7�fˁ��7�|���޵.�ۃVa�ir�K��I/��0�|�_�mS8<�n�ݚ�Н���+�t2��Lq��QF[��f�\%�<4�sg�!�`�(i3�	��x��ݚ�Н���+�t2��Lq��QF[��f�\%�,�F��P��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3@��]V8mbt��]��!�`�(i3�B�+2��;�P����|e"�H�����K��I/N#~8"�Z��l[�Ƶ�1tSjv�!�`�(i3@��( ���M/*�3����3��[<�m��I�՝� s�#���k$ ����l��T���ӄ��!�qg[���**���k� �ԬQ���Kͽ<\��1tSjv�!�`�(i3�o�t����w�`L����Y� ��q�$x=��!�`�(i3i�Q�������=��w)��
=I�^$D���������P�íN=]a��o���H�RtV�^!�`�(i3�<@���ل=����h���}�%Dܭ��}Dq�f�՝� s�#��qX7'��֯���,mk��L�ǀ�:����iW3��O�����%�������&G!�`�(i3�7����������EN.74/���%s����K!�`�(i3�̢k���������P�꠼*d�m�d��-��!duP���2
�M����'����u��r��!�`�(i3h5���=�t���_j���QCH�9#G�>������
�:qEp'{w#/ B!�`�(i3h5���=�t���_j����ۈnp� p��@���!�`�(i3���F��O��ݚ�Н�$f��_Ub����pT�G�&ց�*�
`���n��ݚ�Н�
̛�]���n���G΂�"��ӌ�r!�`�(i3]���\�x8���D�kJe���N�ScM?��y�!�`�(i3�D�������{
Bk	䶙%G�kk�!�`�(i3��jVѭ@!�`�(i3,�˳�*C[��l�,t���H[W?��	P �a��e�D.7�q���f�e�&�U��f�!�`�(i3����&��r��졾�g�Y������y�!�`�(i3�߆�p�h�T���ӄ��!�qg[���**���k� �ԬQ����5��t�1tSjv�!�`�(i3�o�t����w�`L����Y� ��q�$x=��!�`�(i3i�Q�������=��w)��
=b~*��s�������P�íN=]8k��.ͥ�H�RtV�^!�`�(i3�<@���ل=����h�]
���7Ϝ�}Dq�f�՝� s�#��qX7'��֯���,mk��L�ǀ�:����iW3��OEʨ�`N/������&G!�`�(i3�7����������EN.74/�������yr�!�`�(i3�����!�`�(i3�7����������EN.74/���g!�%=F�=!�`�(i3HN��R��bP�63Z�t���%>�rG�@�	������6��+m��o����?c$��!�`�(i3�B�+2��;�P����|e"�H�����K��I/N#~8"�Z��l[�Ƶ�1tSjv�!�`�(i3@��( ���M/*�3����3��[<�m��I�՝� s�#���k$ ����l��T���ӄ��!�qg[���**���k� �ԬQ���Kͽ<\��1tSjv�!�`�(i3�o�t����w�`L����Y� ��q�$x=��!�`�(i3i�Q�������=��w)��
=I�^$D���������P�íN=]a��o���H�RtV�^!�`�(i3�<@���ل=����h���}�%Dܭ��}Dq�f�՝� s�#��qX7'��֯���,mk��L�ǀ�:����iW3��O�����%�������&G!�`�(i3�7����������EN.74/���%s����K!�`�(i3�̢k���������P�꠼*d�m�d��-��!duP���2
�M����'����u��r��!�`�(i3h5���=�t���_j���QCH�9#G�>������
�:qEp'{w#/ B!�`�(i3h5���=�t���_j����ۈnp� p��@���!�`�(i3���F��O��ݚ�Н�$f��_Ub����pT�G�&ց�*�&��j���3��Y$��7����������EN.74/���g!�%=F�=!�`�(i3�U�Z^�t�!�G���-��$�\%e��}Dq�f���4�CD5��E�i�m}6߸��S�Ȍ�kpR,�y6�T�@/�C�1w�R���y+1�����8|��R
�E17�)�#bc�s��HiT˗=߫��I<
���(���Uy��h��G�@�/����t�h�G3�ai��������PX6و�cµ��%��(����e_��|B����$DR�������ן�-�Q�Z�^N�!����;Cj��a�M�{�|Lɟ����I��w�`L�b��K��� �7��a������EN.`H�≶�"ڊ���|��h~���!�`�(i3!�`�(i3p�V�n]�Lq��QF[�b�m��H�\��/1�10�su-�!�`�(i3!�`�(i3?Q�@X>#�ЂDa��(YC-�T^*�h��N�MܻĶ4�Y������EN.�J�,����)L*k������k$ !�`�(i3���D4FF���#���L{����h��N�MܻĶ4�Y������EN.<��{��x� I,���Lq��QF[�b�m��HY'��ݚ�Н�!�`�(i3����oN���[��o}����g�G��0�g�X�q��g��;�!�`�(i3!�`�(i3��b+}y[�Xd��8�(
���||�T^����*�O.�NSG�8�Y=i�&�8nsK������P�꠼*d�m�G�k�a���!�qg�|��'N���+1��y ��/��!�`�(i3!�`�(i3!�`�(i3�_��>νr����e_�WX�iќ����p��&Jhk{��K��I/��
�e~�!�`�(i3!�`�(i3!�`�(i3��'T���+���~=�L���H7��ح4�����o�*H��&��95q��`���φ��<�6�U�7˖�ɳ
xM�v.���)�D��5�v��cg̖UB�nojL]�T!R�ʁ���Mյ���ݑ��3��Y$�M`�K)��v�:�-22�v%��v���ݚ�Н����g!h!����e_�g�+C��sG��Hb� h�ҩι�+�t2��Lq��QF[�Z9�+	�Wsp[��X��=@'ѥ��q�9�ͭ�Ƀ�?PA�g�+C��sc�'�3<
���D�kJ��}Dq�f��	��x��ݚ�Н��H�����K��I/z�
1���;#o�]�ʄ�
%�6W���N�Cٺ��#o�]�ʄ�
%�6W��M*QfY�"Z_�mS8<�n�ݚ�Н���+�t2��Lq��QF[�Z9�+	ҝ'�j
/��ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sJ�A7���ݚ�Н��Ra])n#���{�@֯���,mk��L�ǀ�:����iW3��OEʨ�`N/���:����J0i�,�LD�s�x�-����!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3���M$��2�w����� �.J�>1�Ѯ�a�!�`�(i3�	��x��ݚ�Н���+�t2��Lq��QF[�Z9�+	Ҳ�}�%Dܭ��}Dq�f�!�`�(i3�J�g�*����3���įէ3��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3)�{6�U��(*�O�q�u�PH<!�`�(i3NQw
[��K���!%��v��!�`�(i3�U�Z^�t� "���
w���%��Y�!�`�(i3]���\�x8���D�kJe���N�ScM?��y�!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3:)!�1%�@�	^���yCw�Hm���K��I/y�b�G2!�`�(i3i�Q���'���>;#��Z<��A!>!XM�#����+1�;�.��1���-����!�`�(i3h5���=�t���_j���M}����BK;��t��:!�`�(i3T�=qއ*|X6و�cµ���(A�,"��C&��՝� s�#W���wL�'l/7w|]/(繸P:$�O����K��I/03�� <I��:����iW3��OEʨ�`N/�x{^4��*m!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3:)!�1%�@�	^���yCw�Hm����x�a�t!�`�(i31���~!�`�(i3@v��e��]�Լ�c���J�������n�0R��#���n��*ȑs>!XM�#����+1�;�.��1�>!XM�#�[��l�,t���H[W?M?��y�!�`�(i3����&��r��졾�g��]~ڣ]�<4�sg�!�`�(i3���M$��2�w����� �.J�>�u"����!�`�(i3�߆�p�h�T���ӄb�3�旅Va�ir���J�sy�V��RkB�����X
%�6W���N�Cٺ��#o�]�ʄ�
%�6W����!�qgy�`��vN1tSjv�!�`�(i3�o�t����w�`L���$5� ����:N!�`�(i3C�4M/�Sн3y�ܣ{�j+�j)����r^!�`�(i3��i��:q����J�sy�V��RkB�����X
%�6W���N�Cٺ����J����
%�6W����!�qg�L�[\�"��X� 2!�`�(i3E~X�J��
�M���1F#�֞qduP���2�:
1���Ư����z���B� �b��!�`�(i3�7����������EN.�r6���`�k_�a)!�`�(i3���M$��2�w����� �.J�>�u"����!�`�(i3�߆�p�h�M���yt7�o�*H��& ��0>!XM�#�[��l�,t���H[W?����z����K��I/b�W�
���:�������7�|���޵.��gWaU �IH�RtV�^!�`�(i3�<@���ل=����h�s��m�Eq��lt��T��vR�j�!�`�(i3C�4M/�Sн3y�ܣ{�j+�j)����r^!�`�(i3��i��:q����J�sy�V��RkB�����X
%�6W��b�3�怜gVdxQ,�K��I/��0�|섃Va�ir�K��I/z�
1���;�����u��r��!�`�(i3h5���=�t���_j���M}����BK;��t��:!�`�(i3:)!�1%�@�	^���yCw�Hm���\-{���!�`�(i3�����!�`�(i3�7����������EN.�r6���`������ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sU_GD��W�ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5��6��UH6"����K˖�s���y��lD��~��y8c�D?n����NM���9�O��F����{L,84a��|�&ž_�F��H�����K��I/N#~8"�Z��l[�Ƶ�1tSjv�!�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3i�:`�+PN#~8"�Z�z��B��������p�:��q�՝� s�#��qX7'���q� P�#o�]�ʄ�
%�6W���N�Cٺ��G��Hb� h�ҩι�+�t2��Lq��QF[�Z9�+	�Wsp[��X��=@'ѥ��q�9�ͭ�Ƀ�?PA�g�+C��s���ίݓn�ݚ�Н��̢k�����Tյ���#���n��*ȑs>!XM�#����ևA�d��-��!duP���2
�M���<���H1tSjv�!�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3i�:`�+PN#~8"�Z��mU���p�8���&�Ra])n#���r����;�jmT�#������PLm�<o��w��+-��, ��A�Y�
���3ʩ�E�1�^�
%�6W���N�Cٺ��#o�]�ʄ�
%�6W����!�qgy�`��vN�cN�0*���k� ֯���,Ѳ��=ow_�mS8<�n�ݚ�Н���+�t2��Lq��QF[�Z9�+	ҝ'�j
/��ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sJ�A7���ݚ�Н��Ra])n#]���\�x8�Q:��?��b~*��s���v�)y�Eh�ѮYț{ݮƻ�@duP���2
�M����d��-��!duP���2�:
1���Ư����z����-����!�`�(i3�D�������{
B��e�g�����SY|d!�`�(i3:)!�1%�@�	^���yCw�Hm��!�>!��!�`�(i3�k��^�1�є��g��h�ѮYț{ݮƻ�@duP���2
�M�������xQ�Bvz��Mk�duP���2�:
1���Ư����z��s)l໶�,!�`�(i3q�z����ԬQ���Kͽ<\��*���k� ֯���,mk��L��x{^4��*m!�`�(i3����&��r��졾�g��]~ڣ]h���UZ���ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sJ�A7���ݚ�Н��Ra])n#~x]V�{���>E-�N�&Cd�c��aj�\���7�|���޵.��&���Z����@�f��Lm�<o�̱�	P �a�����=��w)��
=V�Q�� h�ҩ�!�`�(i3@��( ���M/*�3�IX�B��7��q�$�E!�`�(i3!�`�(i3!�`�(i3��D��x0��}Dq�f�!�`�(i3�J�g�*����3���įէ3��}Dq�f�՝� s�#W���wL�'l/7w|]�o
�Z���\(�`���~=�L�.ama�`m�>!XM�#����+1�;�.��1�>!XM�#�[��l�,t���H[W?ð��T�ݚ�Н���+�t2��Lq��QF[�Z9�+	�Wsp[��X��=@'ѥ�!�`�(i3i�:`�+PN#~8"�Z�������!$�8���&�
�:qEp'{w#/ B!�`�(i3h5���=�t���_j���M}����BK;��t��:!�`�(i3:)!�1%�@�	^���yCw�Hm����x�a�t!�`�(i3��Ě�����}Dq�f�HN��R��F F�E̠ʁ���MյK���/C���>e�-�����@:[�Xw�`v@C-�!�`�(i3,�˳�*C�����p���W�,�_sa��o���H�RtV�^����&��r��졾�g��]~ڣ]�,�F��P��}Dq�f����M$��2�w����� �.J�>��2�N�3����ۺ�u��ݚ�Н���w�w:�!�`�(i3��Aڬ&W�����=��w)��
=b~*��s�������P�íN=]b~*��s�������P�ڎC�?�M?��y�!�`�(i3����&��r��졾�g��]~ڣ]�<4�sg�!�`�(i3���M$��2�w����� �.J�>�u"����!�`�(i3�߆�p�h�	T����[
�M����d��-��!duP���2��'��V�Q�� h�ҩ�!�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3C�4M/�Sн3y�ܣ{�j+��x���b�!�`�(i3��jVѭ@!�`�(i3�D�������{
B��e�g�����.ݍ|�!�`�(i3ђw�)�WA�qIp��K/�k�2�n�)�� �g!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok��ʁ���Mյ��M�ԩ&U�)j�S���vo� ��M�#�q9+t�}�ݚ�Н����g!h!����e_�g�+C��sG��Hb� h�ҩι�+�t2��Lq��QF[�Z9�+	�Wsp[��X��=@'ѥ��q�9�ͭ�Ƀ�?PA�g�+C��sc�'�3<
���D�kJ��}Dq�f��	��x��ݚ�Н��H�����K��I/z�
1���;#o�]�ʄ�
%�6W���N�Cٺ��#o�]�ʄ�
%�6W��M*QfY�"Z_�mS8<�n�ݚ�Н���+�t2��Lq��QF[�Z9�+	ҝ'�j
/��ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sJ�A7���ݚ�Н��Ra])n#���{�@֯���,mk��L�ǀ�:����iW3��OEʨ�`N/���:����J0i�,�LD�s�x�-����!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3���M$��2�w����� �.J�>1�Ѯ�a�!�`�(i3�	��x��ݚ�Н���+�t2��Lq��QF[�Z9�+	Ҳ�}�%Dܭ��}Dq�f�!�`�(i3�J�g�*����3���įէ3��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3� ��F�	kwJ�Rmv&&�6,d0����1��eǡ��=֔׹���& d��]�?��\f����ljN5(+Wp��/w1z��ӊH {��u��]'\gWg��	�Z�kfcM��fZ�{y����i�q,?5qօG�j�z q��j�J^�'ž1�|��P�:k& ��-������.J7h�lr�{��|e��0�U+�qbp@�!�`�(i3��$F@S�� 63�镋�%>%���Ra])n#�璓�c�������t �[l;[�G���KlG%��`��ǚ��ظ
��@�U#;�jmT�#��ɂ��.�n�� ��M?��y�!�`�(i3��NƥN��nF���<�W�.�P�	��
�Q�}�	��x��ݚ�Н����3%���v䡩ث�\��N�Ś�-�������y��lD1�7�1 �I����|���"u����O\|�?���-�����H�������U�._���"u����gy岟�91tSjv��V�52SG��E��B�1>3d?���, �I��rʒ	��x��ݚ�Н�a��?p����4��Q� ~��!�`�(i3�5ߧE4��!�`�(i3.�T�+%)�6�Ac�G5�q��e��u��r��!�`�(i3�'�c��(چ���9%����M�!�`�(i31���~!�`�(i3/w1z��ӊE�g�������(ӈ���m�r����!�`�(i3���F��O��ݚ�Н�m�ڨ�hծ!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j�_�Ƭ7~���N�KRuD�*'��>E-�Nb�Sc����E��B�1��e���az6j�"Hs�@�;��@l��O�W]�J��>Y~H<PBn��akaE�,��������!6�o8:4�I���c�90Mj�dL�{y����i�q,?5q}�P�|��U���e��d9=���u��r��J���hB;74/������.ݍ|�̢k���"��w6�0��ɗ��zi#Y)M���Fe��-�����D�������f�\%�;M+�W�˖��_j���?\�z?Xk��;�P�t�5�׹���& d�����9�������ȫ_VBn��ak#����f ȕK�nثIX0F�MV�ҁGG�K�BN
\����+�^n=\f�5>���D�������qD��=a�^7�1tSjv��o�t���>O��T �5�������m�Q��$���͜P_�_S:g�RMm�o��'����u��r����3�Z�#atw�t���%5�����0	�+G�c��Be�A�}�	76�&�� Ӗ�t$�)�vx1x#0<-�1#����f,��ف�ׂ�bƑ�䡺&Y��V����t�T��?E-h���U���e��_	�Ƽ��S�J\7 ��>�:�xjzӝ���w3��׍�&�U��f����M$��2�w������vP8!�>!���k��^�1Aj��t�35L��$
8��2�ֈe1tSjv�C�4M/�Sн3y��'r4�c=A�qIp��K���{#zy�$f��_Ub���uQL+��φ��<�6�pq�� oԔ	^���yK�VSƅ��	^���yحM��1�~Q�4�gX��!z1��,�U��)���Y;e�iK-pm!9�>��n4s1�U��B��-|k������������r$ɓǉ�.y�U=˅ ߛ��u,:g�.XvuD畆J�a$�Y )P<�ܓ�Y��F��[��l�,�nz�����/��kOT�o�t��{��b�b�*k���������|e"������P�]Z�����q9+t�}���������~=�L��i
�i�w)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0Q���
<�,:g�.XvuD畆J�a$�Y ״$(�>g���F��[��l�,�nz������K��I/2f8��E�O`�� \)��\���S)CBg�Xs=ȱ%5�����܋�n焞W���b�0�����C=+f!H�N(�gz��B���=5.B������}Dq�f��K��I/G�?-�Dc�'�3<
�u�����HN��R���ء�I��߸��S�Ȍ o�n�J-\ٿ�6�P��3����!���;oN�	mH����t�T��?E-h��`f���sd�G}%����3f�B7�Q�����A@x8g#��xjzӝ���I(͂��-����^	QW�Q!r�!���;Cw�Hm��K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK�����p�=��d�f4������&G��'T���+ݰM�_�G]�;o�� ��c�'�3<
8����J/�;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�U�0��IuA]C��JJ���L(����7�|V�̹�2�����=�p>�"Y\mJ���hB;��i|�l5R����$~@=7�7K�Phy��te7�i9>���E��xLM[��T�g���bӴ�G�*�K��I/��=����,��	J��I�#�ǖ�޳@�2O��^���+| ����P�D���ׁ{�O��+0◤S%�}t�4\%��t�|v�~�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��q�l���"�aGAZ5h�P��{˒��5��X �צs�6���Sx�#���陋�w��v�9��)�� `l?��f��/_�J����B�����HN��tOIkV�g�uu�i��b���nu��3�����-!�ρ�G����8�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�7_�|{�����X�혨5�����h^���s��$�Z;��|B>&k>�Wz;��|B�I�����
�w�u���	��-���](ùy�;quA0�e]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7���_J��`�k<�*y�$\���F�`yx�>�+X�[�G���K�k��M����$A���A��S/��kOT�>���Dl��ִ���	ɩ���@|����^a�nu4Bޗ��jw�	���@��v{�G��R:k�ڛ��¦��ѱ�R:k�ڛQF����㔐�H/��fm`&�[���a��o�����]�KS�pT/�GS�⽥�R���h�?�m}}�G�hA�3!g��ݚ�Н��>���Dl��и|��?�Օ�R\��>�������Ra])n#���r�����d�tu�z���?T��'�PD�HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}�-��cR�O�������Ёg�#
VҶ���T䤌ZN����6�o8:4�I���c�90D�O�,e���`���φ��<�6�^���+| �p�8?�e �H����Qw�c4~Nr_�mS8<�n)�{6�U��eX�LG�5:W�^�|��/��kOT���=7�ŷ�{z�n)P<�ܓ�Y�߆�p�h��d��JXl'�T��~��?u��C@�ݚ�Н��G�-!�5/�V�q2�Va�ir[��l�,1B��CSkG��Hb� h�ҩΦ��=7�ŏ�ʳ�(�)P<�ܓ�Y!�`�(i3֒���\��#QSU:�����|e"pT/�GS�x�� U|��v��ONH!�`�(i3E����[����>^17��"��ӌ�r
�:qEp�;�P�t�5!�`�(i3����/��oځ��p��^"4/����hu�A�">u��r�幁+�t2�4\%��tF�̃��H��}Dq�f�$f��_Ub�F�S�1 ���Ě���fR��}���;�P�t�5�Fr��jZ����~jܶ���T䤌���7�Y�(�JZ�Vk�;��|B9B�X�.o���C��m;#��Hۭ/!�X���XXj��9^�cs�C�(4&Ƒ:2�c<�^<�H�;�pY�Y�|�8�ܬS-l�ݫ&�b%%�Jם��S>������3'�2�@`u:j1�e�Ǧ�Mj�(ȅ���2��.�g3Zv���� Й��B䧹�$�=�}!�`�(i3!�`�(i3!�`�(i3U-��_M?g���Οy�<.��2-@`u:j1�e�ǦU��֜��3#D�<�O[֒���\��x���"7�΁M�$��ښܔ??Vi� �Z�( �B��6��#�?�B�b���ߑg�Dp��H�ϋ�LΗO!�`�(i3@`u:j1�e�Ǧ�5�%]���a(􆿳�ټ*w2�564��X:��K�
�M�J�g�*���p�xbE�@�̔A�qIp��K�s���.(f�L�#�E�fD�GB<x ZR��p��ύf>�Ns_>5m�,�D�⅒������q}&@��&�����	��_$ر���闝��Ν3�x���(hyX�[Ӿ�h⧂=�����ny��^�<���%� �S3�
T7#��ג�$�3��4c�x#�}��6�Rh�HLN���R�lD�GB<x�o����U��8��6��{)i!r@".M��lqꨳ��5����`Kn���P���Gg�R|��'=i��)J��P>�%��v��Bn��akl��X|P����t�T��4c�� �܋�n焞�v��A)��Ҷ����S��R&.'/D�&�8nsK��\���S)�K�U���;������tD�#k0����+�^n=\f�5>�1x#0<-�1���%����Fg�U�D5�v��cg;�������8���Q/�"����,�[��*c�Ѥ����vo��VF�˷��%5������Ҷ����S���|�a�\37+�p�����U^�Mi~_�T;�jmT�#��\���S)G�6�!~�#o�]�ʄ��.�L�oDy����ҡ"#�k�	���QC�0q�#��d9=���u��r�婽��&�� ��\�&ɖ��_j���B~?X:0�C�l�kZ�[�[]�M��L��}Dq�f��k��^�1g�G��0��'���C&b~*��s�/$�ߺ��]��pZ�ì�d��-��!g��J�s��{��b�b�*������� h�ҩΖ7������8R ���M/*�3�2�:�#LAY���&Y'���4-Y���Ra])n#����,��=7�7K�P�l[�Ƶ�	���QC�Ҷ����S���Cu�;�R��3��m���d������z����-����!�`�(i3�,�B���{
Biۧ˺�s�˭;{o�Ϧ����ھ	!�`�(i31���~��+�t2�;�������w�`L� 1�Z����o w&�s���%>�rGO�D mWNG�&ց�*�s��������2�(��w+?i�Ct!�`�(i3���$A�;�P����|e" ���Aؠem���d�e���N�Sc&�U��f�!�`�(i3��3�Z�#aȮ۔��5��Y��x�1�-Ϩ�ݚ�Н���jVѭ@!�`�(i3�,�B���{
Biۧ˺�s�˭;{o��n�(Z�ɽ��:^E��HN��R��bP�63Z�tx6@��� ��˭;{o���XW�G�<���>e}I�6������U5C��r��&�����&G!�`�(i3U�07�:�tMɶ���74/����G🕾{!�`�(i3)Յ�N���^�v�����;q�"��ӌ�r՝� s�#���k$ �7������8R ���M/*�3�2�:�#LAY���&Y'���4-Y��9�O��F���R:k�ڛ)�{� �"k���������|e"$f��_Ub�F�S�1 ���O���b�z'hۉ)��ipɳ4?�{�XԔ�Z?�߸��S�Ȍ^��,P�H�*U��;�P�
e�,��P�܅��+jq�����Å��������lz���AZ���d���!i���8-|�D�"Q�8��߹�q^�j3eD���w��=�Б�����ph�)�w|�0)��]��.e�����م���R�n_�A޿b�i9������ћ�<�����k����=��ʊ�z�]���,��"�k�;{���Κyfx���f�Y�����M�!��^��Bc�"�"��������k����=���_u� Ф��,��"�$�r�9J��:������èVp��E|��c�S�u. �����n_�����S���� "5�]��'T���+�Zn��޳Q�4�gX����cl�"��Z�Z!�`�(i3��w]��&�4>��K�&Z0Q���s��5�q	��F{/�����,([�y�
%�ǹ>O�-����`����줞�l]��SFU� �h��@�hGq6��nX��U�	vn����R�����_���!�`�(i3#B��F�!�`�(i3!�`�(i3��*�{6�����&!��ȁ��;�<n�f}�T�NHX��+���;���5��K��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3E3����.��FO�&�r����'��,#�@�΁�a�n���X;p`��vbëdP3z%�u�܆X:��+��b��v�#$�q�
k-���w�E�V{�!�`�(i3?�ᒹ�G�!�`�(i3!�`�(i3���BjJ�l��!G���r������z�r{]i!�`�(i3�X;p`�U��֜��3��e�E#��!��B�R��0����ݚ�Н���*dy�ZB؋�Ly�H!�`�(i3�P�Kf�h���J	�J�y��*?(��N�����~Y}J��F!��&t�ND�����X;p`�T���'/�>X�o|3�D�c�J�.��8z�f�h�\ƙkH*W��u�a�ݚ�Н� ��ߕ!�`�(i3!�`�(i3k S���z A����;���C#����d�E����'m�|g�~p!ۓ�ݚ�Н�&�2�������ȍry��	��b~y� ��&8�,��Om�"���^��r�VU���l����S4�0 L?�p���@Z����
� �!�`�(i3B��亁���&�%���B�'��a�[<�!��Tl�������l6��Q9���ۗ&8�,�cop ���6�G|��2��}����a#�fS��I���i9>���Ef�?ǉ�=�e�MW���^�yO�j���H�D���dݮ%*!�`�(i3���_͏���/ӳx��d��]�Q��f�_���u����g�&�0m����#oMS����6s
�:qEp0���Y$�8�$��`��7dh�?8X�˞�DG�e�MW��T��b9���ey�E�����$���f�?ǉ�=�#�m�-��Vi� �Znj��TAn�OZ@��5�h�ʪ%��18�$��`��UB�L5wG�!�`�(i3�:5A��p]M�|jHX{�t����՜�%P^���H> ��9�/�q#a�_�`�ю��x�T��ۇ�Qv�)�ˌ��Pg<\uu�����r����!�`�(i3!�`�(i3!�`�(i3�z_n�ԁi ���=��?�d���&���d.q��	����Y�!�`�(i3!�`�(i3!�`�(i3�mJ�0�6��"Q�8���������9P�Y�/*<!�F��66����~ω(�$V�y�2�x�h������M�!�y:i������M��j �M1����JV��GB%p�  �fAany�h�t��4����)\=��A���i9���Qp�	d��2������<�bሻ�״:��JV��GB%p�  �fAao�F)���;4����)\�uv�>u��d���!i!�`�(i3!�`�(i3!�`�(i3Y��-�ݼ�յ[+8�a�)��Ƃ~6T���Q�x1�~g_�,\ަ�It��+g[�Zt%��m&<>��%��JU�a�(�n����62�tϛA^��'T���+M�Mb�:u�w�vG�q�:�&����#|�1�0j��*������Э~���V��2
L.�X;p`��vbëdP�4e���>�f�?ǉ�=�1_�
774\51�]2�t��MJT��
!�7�R�"�*}#2\z��``�ǆ�!�`�(i3�&8�,�aG�	�AS3f���])ܟ�Ma`_��r����N�i-9�}�~���lscX{�X!,!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�;�
Ơ�*�6�M)w6(��.�����gRI/!�`�(i3�Y�M����4Wt#��5Z���r����ؾ<k�[��x�ܽ���X;p`�T���'/�>#2\z���&�3Z�K�!�`�(i3�&8�,��y��ЉT�9e��/�7�(��.��?�!�`�(i3t$Q���V�T_��p�V;�������gL�4�2s��2 !�`�(i3��5@~JuM�D���!�`�(i3W�4�:*n~�<�&��Xh�hk��a��OY�P�CQ��Bރ;�{��C�{����K�7��(�mWƒ�a�}�$Ϩ�;?���*/�|�-���w�E�V{�!�`�(i3�;���5!�`�(i3!�`�(i3}���/+��!�`�(i3M�&�mU�w�������*����	�?h���5��қDO,\ͨ܉p����O,8�ݚ�Н�7�N��X;p`����$AA�:JϮ�MQNv�2!�`�(i3�˺�Q���f�?ǉ�=�*46;�[-��$ϙRl�bu�	?�cx�Y��j3����(�a��>N0Θ��ݚ�Н��0V32;5��X;p`��B�+2�A�:JϮq�\E��0!�`�(i3�$�~c/�;���%!�`�(i3�#�l+G�)#��(ߖ�3E M0���M��s,�?�k�V�?�҄���>�S��I�����T7��v��w�K���&v�`�Ll[,�)Վ�a(􆿳�E��-�*���ߠ����9
4�٩czZ����N��E�Es���Fz���w]��&��)��>.$5<�`A��_iN��E�Es!�`�(i3)�{� �"��/ӳxI�؉P���Of�`@T:j�v�!�`�(i3czZ�����oͷ�����ǖ�!�]m�(�h@)í�_�ߍj�������� 63��p�@OM.Irv�-���w:�4Rʹs=���|�F�x
lw߲�=O��{Rv�f�A
i�eL!�`�(i3!�`�(i3!�`�(i3{�d"����MjئO܅.�g3ZQ�ͼ���ݑ/ٝ�r)�!4�,*�!�!�`�(i3!�`�(i3!�`�(i3��/z*q+6j�"Hs�"iJ�����E�a2j�Ph������m�\cw��TN\;�6
�P��#��s�'	�?��[n8�A�A�I��'���I�Ūe�M������'n�^0o��t��>ea���]n�� V���	�e��`������/�_�/�h3bU����P�5��t�l���G���e`Ez#j���8-|�D��*CTR��˹�'O�N+��T��Rc1"�>_�q��.���:��)gi����S���� "5�]ޥ0D���3A�)Oq�i�-}�[�����U4 :��	��aJ �!,P�H@��&-���xԞ�����i��E����p��x.�Knq,���9^-���2��̪U��֜��3�&8�,�e*���	&���`"�G����?�s!�6]��E[WͶ
�`��~mi�ݚ�Н�EfVNN�0|]<w:��X;p`�U9����u���q����k��,��C:���2��}��=�lx+~�S��I���i9>���Ef�?ǉ�=�� ߌ��-��Vi� �Z�xOQ��B�'��a���p��b����z1]�xv�:��p=�n�Ԓ��K�u�c�$�~c/���F�ƻ!�`�(i3~n���,a��/ӳx���{L,8gf�mk���b~y� ��&8�,��Om�"���^���F{/�����,([�y���㋞9�nX�8j
Jt��)���l\�6�'����7Z��$�~c/~�O�������+�t2��ӱ}�tMTl�����)��.��f�?ǉ�=�M�g����-����b=��y��j��k�lԇ�-{�4�0 L?�p���@Z�6[��u�V�<�nbBIճ��)��]m�(�h@)í�_�ߍj�������� 63��p�@OM.IrP"G�wk��jr�!�������,\������,Y�I��/^�=O{Ue��*�̞��>��vbëdP�D�R��	ܷ�4D�P���I`���jVѭ@!�`�(i3!�`�(i3!�`�(i3��7I���
�)W8��V��	��y�㘞������8I��2�HF�M]y��Z�/�N���N
k��L����4��>���O6�o8:4�I���c�90Mj�dL�{y����i�q,?5q��N��)�Q��l�'ž1�|��P�:k& ��-�����D������"r�V�)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b�Ж7�����5*A�u�������$~@l����*��"���l<o�;)�y���ƚ_��}�	76�&�� Ӗ�t$�)�vx.F<!W���zՇK����3Ah	)ޟ-�b�+�