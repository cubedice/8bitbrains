��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�S�T�;Ϗk[�^��_*z�w4G� ������[���a�8%`��4�s�6�XAoeu��a@����þ�V�E`Ԏ��%��1��*�"��Yk"1/���%	v3����M7\F���r��C>C�݂�N$��/���	�0���'v6�o�"c����A�&�8d�v��x�۔7�D��:�b�#�Bn	����I@beB��H��>I��4��u"%�������j)j*[��HMi.��>��'��E����F�A�y]M���y�.!/�1 T�V	�tL��	�<�A�}Q�� �P�_ߠxR�	�$F5��wx0�<����O4��X��m�� N�X1јds£����&��ea�8���*���g S�7���I�N<��;���u��w)�S����w�~篟|�Zl�~�4�,���$'8o9����E��lU��l�����開��g_���L��׹+�o P���t�	�1��"w��N�˥���\�4�sP	�b\qB����U�7��W/�He��ɳ����~�MUs �.Eٓ�9�:�T��|��=o����"���	x]���Ec��$�~篟|��~ ����1�����8�:r&@K,s�θ�<�"������p<�������,�\gE�y�7��������Ψ�w�Ua�21�*��ϕ��RL�a)ѻtUWR�N	:.���n��R��̺~�v#�,�}�7C��H�����"|�Ћ�i#�t{�Tl8��`e�TS��\�4�sR���i1������"^Y怄&��b��~�MUs a"�x���2@�+���c�#s�0���!Z:���:r�a�u�����!�M��ED�D ���
r:�����u��w)�SU��T�d�7��Mv�9�E���5�n�ﰑ��m18�:r&@1�+Q�<Ǵoe� 2m�!=�y����h�}
�ԟ�d�fY�?hP�+*�D^o?�M��;]PF�$8������D҂��9���1�E��p��qx����-&���#��*ά�1�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc*c5A|�Y^ɚ�Ȗ}��*e�q�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ���AOge�Ѡo���h�k2�$�����(����5�2���[@%����nEA�X�f8�A����Y�{'%s�5o�cf�W+`�x�oP��@t��4�u>Kw����qc�U_�+X�p^'�&�Z鎬�����ת���A��%���׈�Qq�Mݩ`~���H�=%+]Bo�A;h�F�`�"Q���]�!��s�XZ8E@��{��&�k�1 �O�oc_����+#��.X���*"v%)��Qcm h��\�vņ���s�c�����gvEU1��?�"��J���T-a�ؕJ���˿��2=+��׌#�����uTo�_���
.���j"�E�	ZE�M�@ϱP}��O�����:�����開`Ai��n�N�Q9���mj]h�E�!	�J�%�XB�&�=T-a�ؕJ�9�#=�8%T-a�ؕJ�>�5�0���6C�&/����D�����0�$i��k�eǎd .8��|K�{ߝ�Fc��B�I%ji�7��
#>:��� �rmd�&l�����i�I��M�3q��=$���A���ۖ?3�'����1Y�ΊS&nQ�rV�kV�џ�}$|~ïSup�xg���m��T���u�Ia�6~n!5�$��fP�_�oK��͏x�e�]�c������uRBO ^�̒��b�|t���o�[�iu>�$fwa�m�f�#zX�����N�0�/<�U��=>bMM`)��5i׈�1^��W��E��e߃����XRe><��B9'���Xw՚�છ����a�"Z鎬������	c�u���E��e߃����XR�[R*$�s�,�TMo������a�"Z鎬����:��q�_�Ã9���1�+��T����oGo�Z�J��ݪ�b��颥��3�7DY��S�\6��L�͒1�:�Ω�S�T�;Ϗk[�^��_�9���$1me��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��ly�(&�N�����B���0o����T/{$m)mW�/��)�-��DǷe��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�I�+�c��Uwz�@ʶ��辐�!JHn��z��C��ྐܼ�\�v�9�#=�8%�b9���J���z�my±�sR�{F  M��va�{����PD}#��ůN}�m��{B���T�D��\�v��8&���I���8|�L�*�g�;�k	�oG�� h�ҩΣ��n����-�����y��j��k\y[P޽��5 cd��#�xy}�����H4 3g�Y�T�:5A��p��jVѭ@�y��j��k\y[P޽��5 cd��#�xy}�����H4���b�%3�;b�-�2��;�P�t�5��w�w:�;�jmT�#q�P�:땗� h�ҩ�p��xs�S�*
�DWo$ۯ}z�| �8b�9A�i���Y-]�\^M�Ɣ�	��x��ݚ�Н�
ҭ�3���#���1��t�Q�n�!�&}Ji��6���l]�a��}Dq�f��5ߧE4��HN��R��bP�63Z�t�y�"�V��5M��z�o�*� '�!�J����ϩ�Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����m2����H�� ӫ/��m�Wq�
Z*�)�J[x�*��rC3�8�c㚂�IB�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a%��b����xVg�uP.},d�z�m�~�.4g$�co�XB�&�=�b9����N��a'��@��(5-ˤ���k�˒�����j�'l���u��-���E�0w�m��<�mlo�2N��n�=U���iAe��Y��)�?Z����JHn��z��x�f7﹏,���D��a�si՝ӣg{��aDeq��ҝ�r<�n"��g�LX�,T ��b�FP&���rS�h!�`�(i3�@��O���Қp%�0�ΩyO^~��M����A�m�(��ڽQ����2N��n��t�J�Yy,P�aw=��E����F�_����ֱ�q��w�G�ïWA],S����|:��ͼ�\�v��8&���I���8|�L�*�g�;�k	�oG�� h�ҩ���D�Ώ�ƅP�!�Sbb�����@|����r�����L�����U�ჴs3���l�c�5ߧE4��$�[��= -|�GP���*y}e��p��G]@w���a��G~�= cZ�-ڷH�%����@|����r����~Ps�Й���a+Q�� ��s�gJM!�1�� HN��R��F F�E̠�i7N�_�z*K��I4��欱���j���]���.��|#HK���v����`!�;��!A2�WA],S��o1s)�u��r��o|���P��3��/���WA],S������=�՝� s�#���k$ �<�I��y�fe����~éޝE��Qfĉ>99��A0ok����DFTޱ}b�g3�UX��xϚӬ�5n��/0�E�i�m}640�RS���$
�)N܉}�B>i�a�	KX\�B� �b��֭�h��O�Q��ǺΕ�A�m�(�O�Ŝr{= { _Ta�F��l���)�4�����Ὡz�*<�����s~��!��jVѭ@o|���P��f�Nd+l�Yҽ֗��Ǒ�o���D�Ώ��V�:�R�;�P�t�5�37y�����:����@��%/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!�_S�t�Aju���lWg����ha�`�2G]�Mq�}��,+$\�M���5E�[�c}�sX�>P�2-i_�	,JZ�!�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�NilM"�����iM0�3m�:3��Տ�L� $�3"���N�T<1(�d���Mo�~$5��_������"~6���aq�����4�k�߻P`���;���N���M��A���va�{����2����%��/q|��h�ӵeoQm�`aĉRW�F��F�zL͊�q���Z����p��J(1�:�>�̸��oJ(�c�-1F�]�q:��c^�Զ]܆�����ң;�f����~����y�Zk��~��6n�L�%��/q|��fx'v�ao.\C�k�Ԝ�6NzL͊�q��]� ���_�hbvk~�#xB).V44�o�.ᬵy��ՙ�3Ќ�L:(�
�*S|ò���
��_�����k�79�����\�v�%�M�5&l����I{6���>�3���/��¬3T���&|���BY��l��=5;���ip>��<ug	h<��Q�R{�lp�q04?VS�����ud��%BJ�g
�zP�w:Ec�[�p(	��Q�^�y�zL͊�q��j.��?�Uʚ7�ܩ�.fOe	�o1�ֵ@�3���/��;L�=Q ��b�FP&����҅JHn��z��`�+]���e���im��mų��n��Uʚ7�ܩ�.fOe	�Ƞ�d�P_�n�To�[�}�~��l�}`V�u�6������1�R+-h]��.�{+�&f��w�'�4uB���u�~����J*�Rs�0K=X���d��J>�߯�"5�o٥����Y�JM�b��v݋N�����7u7҃Q*�6������1�R+-h]�83NI�����w/,g{Y#0����l��=5; �e�B�R���>_�4uB���u�~����J*�Rs�0K=X���d���fx'v�ao.\C�k��|��-�Vc�$J�{�����~�=��K�I0���ԏ�.fOe	����4�l�>z�Vg.N������[� �I�������m��b��v݋N��������џH�5ߧE4��?"�����2$%-����y�����=u~Ei�"2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE�7�0}7��k+�=Qj#`�,�mI�p��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�Ia�6~n!5�$��fP����E"�T��b9���M��A���D]�$���k�1 �O�o/��T�n*�N}�m��{B���T�D��Ψ��F$��O�&���e�JP2Ud̞��>�1���t�<���8-|�DOYZ8�%QQ�{��x/��Qu���%<i�LE� R1Xi��&\})����K����J���y��j��kj�����N�_9�R�5;�Щ�j#/M��\�jX��u��A�0�Ή*��a��Ɇ%5�����{��ü��O��b��֔N���c.�'}-�����@E��=�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��0���V��C�qҢ�����N[ m�N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開�Њהt�ȳh�L>sP"G�wk��a�S.l"�S�)37J*u�1��r�p?��$�Qu�&�<��G��d�٣�����c����յ[+8�
ҭ�3���/��kOT�i7N�_	�z�w.{��w�_��(�6k�4d�{j����·/ҳ�ϾQY�u��A�0���򴶽!�y�"�V��5M��z�o�>��U^[U�7�tW-�J4p'�>��\��:��Z鎬�������(���w�?�b�>��]�!��=���W�N}�m��{B���T�D�]�!��`��j(&�L�i��ko�$ƍ2���lĦR'cf����T�x��QU���^4��y��j��kL1���oB�T���I�!�w(�y?�?�JY�)�֬w�J%�H���3�}@��9�ڮW];��e�8<�V�Zs˿�}w��ea�8���*���g S�7���I侰j���