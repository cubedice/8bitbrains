��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}"6�l�:���L|�w.j��6��H4ي��2_)��:B!�b�ؐ:�{T�{df;���a,xh'�$k�w�D1���}����ň���x�w�Y��k��ı���$��������j��t�w`ۺ����N<��;��� B]�pE���	x]̃Dj#^Da����M�$����o��I�绯�t�z����)�,�˛D��w���旴4w�1����h���������$[Z�i��%A�a��gs|�e
�9��Ax!P����9SA��R����.���Zߧl4���0�?�1~�x�c�� ���"����j�͚L�	
o�;�i�8>'f(l����x��5�O���}@��r���7Ȭ�ϏI �ol[�y���Q\�_q_�'�i���m�}�Ć�,I�@�"|��Ca2�]вk0��}9)�Myիnň��h����c$����k��[/��ԅ1Qr������i���'d���C�0�%��w�Q�r�4����8ZJ*����	��ZHz��	�zy���i�!�`�(i3!�`�(i3!�`�(i3,-)��8�g��F�蹕�ڐ6|Zk/�/�}���1�1�ҕ�/37���E�D��`X��$D@P��f-�*��IHYH��cJė/�Ҏ�|O���4d!�`�(i3!�`�(i3!�`�(i3ɬc��WNPw-�h��� ��,/�J2���ں��)��'��8�-Zy?X��/4肋�FS�0���>E�C6?6�=B���:(̜����,-:���h�;+3�&�K5A�14P8�!�`�(i3!�`�(i3�0�9&،EB���w�[T�� TY�Iݹ�ˀ:��n�7�����O��t�sȸ�"rR!�`�(i3!�`�(i3R�����Uq9�w��Yw߿���̙	,N�Eĳ-�)�.|��]|F������sȸ�"rR!�`�(i3!�`�(i3��,�0	C}!&��[ܳ�G���������{7$0~'��&\VI`,�ʺ�;[��+$�6ﳌl��t�1��꧄�c����E�zy�զ3�0�jT ���#J��;R�S�!�`�(i3!�`�(i3!�`�(i3 ?[n�:#G٪�t6�yG�?� }[�KO[2vj���B�N� ��b�FP&ׇӭ��!�`�(i3!�`�(i30R��=�El����W\0���JY���y�!��_��0�/ᜒCX��)��h��ׇӭ��!�`�(i3!�`�(i3I����CWI�R��R���w`q��&\VI`,�$��*�z,|ފ������o������$�@�8��ˮ�ڠ��N�[�K5�����z1F~�����8h�M���W� g�[�ܣ(O#�e!�`�(i3!�`�(i3!�`�(i3�y��ă/W��G���������v��_�f�z�H�}tގ:��sȸ�"rR!�`�(i3!�`�(i3���ׂo�4�)�y��L�Di������<�FxNߡ�����Fz�!�`�(i3!�`�(i3�H�"k�j�EB����
'��(�<&���@��� 3�
2��k�B�p��mAe�sȸ�"rR!�`�(i3!�`�(i3��؆�}X�6���j\�d��'��_�]�0��zO�)�C�o8�����i��1�x����NQ[��Y���x�la��jPG���7���6�!�`�(i3!�`�(i3!�`�(i3u�+��{� ?[n�:#G}��F%���B$����&\VI`,�=JK�t���Z.�\�ػ�G�E@��j�g��o��/\k�l��p!!v*!��G�$U����ߪM3��)CSa��KlgI���7�����3m@!�`�(i3!�`�(i3��+�t2�8���]���[
y�s��;g�(ñЍBN��ç�"$�3�}����Fz�!�`�(i3!�`�(i3��p�!-�8}�����'��_�]��_��05�q��e�Ƃ�];/��������Fz�!�`�(i3!�`�(i3�*"�˪T��$�} ,`&�}�؝�T���ܜ?n昼�2#:�ֵ*&E�^8��xt��:_/�~8����A�߲wb��� ��WM�P[����(,)�=!�`�(i3!�`�(i3�B�'��a�{�ç�o�����0����(R\֎u��� Sgȼ�sʫ|H�ͩ�QϿ�ey��<0!�`�(i3!�`�(i3!�`�(i3��sƲ����e:��x���ᐜ����!���C�/�y9.Y'`f�������
��H�ƈQ�H��ޝ���'QԤ�7���6�!�`�(i3!�`�(i3!�`�(i3�7>�����D/͘B�5�35�#� "�q=i�/�J�0�)�u',�G!�`�(i3!�`�(i3�2 /��u��
���ƸtU�����*��>i�!����n,��'�\�n�~��q"P�H�oe��C��c�S+d�J�Г��f�u�����!$檦!�*��Q�`��=vݖ6�F!�`�(i3!�`�(i3��7���,�K�!5�����n,��'�\�n���t�u�?9Pjp��h���~�I��J#�2o�lS��?ꆂ�5�80�[X�b\g���J��<�i��o�]�E�%X(R�6���G<�ok��u4�w��dr��l"�X[{�25�M�1�>�J8�����È���_����Г?����."���T��� ���8ZJ*�`��Ā�	���8�� �Ļ�Q�?���c�r���q�sϻƫ}�=�������d=���q"_�v���Š~r��<Y�d��Z���붋"�M~�7>�����D/͘B�ۭ؜�J��Jt:��v{t��qS�j�e����������,[$��.`.{Xan:�ke�"�q=i%ʴ�ɒ�L��C�/�y|2I��js�B ���Wʂ҅��g�������������(��K.����M
�a��A@�r$��k���:�nj������y;�j���F���+2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE���Q��f�SR�v�����������\��o�?�m݆�8m�4|/yl}Vİ�6��$�.��Ԫ^��rL�%�7��Ŀ<Ԫ^��rL��c5����L�^
��r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!M�c�0�gB�1���i�D��0�������"��g_LG4A��/���N9D<���]ȟ!�� 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������ݧu7Y�M�+|�#��Byl}Vİ�8�d��N��yl}Vİ��8m�4|/yl}Vİ�6��$�.��yl}Vİ���Q��S
�yl}Vİ�M�W9�f^�yl}Vİ�����k0e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���2O��'HY-w�Y��k��ı���$��������j��t�w`ۺ����N<��;���u��w)�S-!������~篟|��*�A���I�n����fџ�_�v%�~G�6֍�r`_��*�u��.t�5�M�1�>�8B���<{��*b.[P�x��t*�=�V��u�/��m��@��V��=B��,����t_Ȥ�W�w��fD ��b�FP& ?[n�:#G(+F�	BaN恔� 90'�f����&�&�
.�n��������SiC���\#�t�����ڕ�>���??[�o��RL�a)'r�Ӟh� mߍu�M9�ߤ����Q���@m��7C��H!�������0�'+��h��=o����"���	x]�"�PL�,eHc�J�M=���-�:1,ĠԜџ�_�v%�_ y�+�3F��m1G:��"w[&�K!�#n��]t�#K�{�:H7ǫ�V���V�/)�Myիnň��h���|~�@����k�8���҆�|n��)8P�d'�%��hݜ�����AQ6|U��<d�L\�Յ�B�U�٣�R��$���"HX��+��^gg1�
հ��C��iF&�A��h������:��KL�����.jB��@۩�����k�8���҆�|n���&�]�68��hݜ��  Y0�����N��%L\�Յ�B�U�٣�R��$���"HX��+��^gg1�
հ��C��iF&�A��h������:��KL�����.jB��@۩�����k�8���҆�|n���h��C d��hݜ�����aj)�>�,r�F@�4%������I�Z�*�I���Ϊz�&���Ḱ��fM���v#n�0؈sU����A����&D��0H����RL�a)ѻtUWR���I����gy3�]	��>	|!�zg�Z�$m�a�gPM��r9t���k�8���҆�|n����{y�ڗ�B�����[AF��ѕ���<l���9��Q��CpC���D�v�{���c�5��<�>�N��̴�*V��z,L���	x]̍��;������#x��(��[�� +u��Ix���y+�����S��&h���y���La��;���g�Ȝ��@�r�O��C��0��$�>��w�*��D����Ǳ����w�>��SX`X�B%�r���7ȓC�-`�e�g��!��x���� �"!B�������.�-���
E�HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�
+&�s�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�f<�,=K�F�~�����J&�������[�/~/�ח۲�J�[j�fTܷ��WL�C�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ���AOge���wV���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcC��M%'.V&��B֥/~.)��3\�R�F*}�c}��uO��������	́߶`(r�M$�*�X�f8艢��S��������Ǜ岦�%I^��������D	��U�e�n�^��]��g3������ɤ|pW�Cy�w=�4e=��-��ؽ7$�	�s}��[�wH�HͶ���ܜ?n昼�2#:��b9���P9b��	�Y���1��� �U��֜��3JHn��z�C�$��؍��R��j�.(Wx*�_F�k-�!�`�(i3��|g�Y�'���Xw�������펎��{5Yl���#��]���>����Cί0C��؆Q>�[G�-X�@�^��1�(R\֎u���sRt�7G#+��\w��0](@X~�H:�W��7=c��Et��q���U�[��N���v�Z�]2�y�Z鎬�����	�7 �#�\1^O��0ˋ��I��w��,>����C��(R\֎u��ԟ'�D�7G#+�Ǘ0z�cULy`�_I�v��4���OTWRdr�Jbk-����'�\�n�wa��>���g��U-�e�,���6+�=�B4˖ב����E��@IE�U��*�QN��� ]���f�fx��V$�w�I�?g�f���\X�<����8��UWJ��)��q鋴�*Х�]��:N��;
�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h}|��XH��9��p#�7ڜ¸<�X��/~.)��3\�R�F*}�c}��uO��������	́߶`(r�M$�*�X�f8�b!��u፧���0��G匵��:
��]�!����w�Հ�(.V����+��\��ޡ.pz�Lۘq���U��@����gG=%� g�Vv���y��7s�9���o>��l%i�-����]��O�M:R	�G�L3cfi����hD�v�l�Ū�TD���)T&I2WM�vT�V��|�������c�A�L'��~�2�?�B���N�gl��ܬa(􆿳���2����.��DP֞ E2�DZ���ǘ�g��O�M:R	�q�W:�m�N>�4�
��S�,�:苙_���<	�Y�{'%s-�,�c��g����R5Xx�w�?�b�>��]�!��	Ǹ�y85����XP��~�26��\�eK&��s��a�\�����fZ���o ��b�FP&����҅�d�٣��c�A�L'��~�2�?�B���з��H��g��U-�e�,���6+� ��b�FP&�%k�����d�٣��c�A�L'd���v��R�wX��d=��¾ȼ5�����}Y�5�{4\��ƽ!61��aUp�rP��O���2�!�x=�FZ���7'��U�RmN�sA��6��-�˫�_Q�D�mu�e���PO�my$�N��o�/���;��6��X36$��&�D�muշ!Rq4������!|P��ݓ�W���KU}>�<zݠ�m��/�
cFI_[f����It�ʁ���Mյ���(��L?��:�wǹ](Uy��C&��G�&ց�*���c�13�h�6�q��S��L�e[�8���&�(*�O�q#q�;?���2N�3u���Ǥ�ܜ�}Dq�f��x����ն�l�P��j�/T�<�_˻Z�}�ݚ�Н���5����@���Z���{�u1H3�AP}܊�ti!�`�(i3[��4��IR��������$t���'i��������6��u��DH�q'�D�mu�#��bE������!|P��ݓ�W���#
/3D�rݠ�m��/�p�c�Zf����It�ʁ���Mյ�$�㚬�L?��:���7�3m��C&��G�&ց�*撠���\�h�6�q��׈��}\I�8���&�(*�O�q4����T�p��2N�3u�gl��̲��}Dq�f��x�����Cv�#!�j�/T�<�_����/���ݚ�Н�)@9� ����Z���{�u1H3� �i�7�*!�`�(i3� ��F�`���A�P�$t����ıA�W�fĉ>99��|��3��H����	�44�38�Z��\_���ľJUp�rP��O��F`S/��7>�����ǚr��y�!�W�&F[!�`�(i3l��`]*(�I���w�:?{CW:�+scX{�X!,N��e�� !�`�(i3!�`�(i3!�`�(i3rW�F����Q����Y�=�BZo�7>�����ǚr��yݥ��P];�֭�h��O�c�seR�a?��`��yy�RA<,�l�}�L@t�"�5��.,0=]^	�&|#9���Ra])n#���r�������f�R�{y�Jܹ^�V]��}��Gr����L��R���}Dq�f��5ߧE4��HN��R���מu��� �H�0��
�y�"�V����譬��f���,9�h@Zd\a�U4�1i�7�cL���	Ǹ�y85���w�%s�iI9�o�L~΄gO�3��|��[��5��S	JZu`Ʒ%k���}o�@EZ����<Z��u�=:�NI+����	h��4��+��\��բ,)1l",oMG~�K�3�Ƅ�u",oMG~�v��H���������%���h� ɤ���ms��/�u���4���O�>�k}�r�����Uh1�;��|B\�2�R�G��%��ڽk�5,���������9b�S� 7�v�ԯȥ�����S�7>�����ǚr��y�#�ϲ XO�M:R	��P��<r���;_��8W�w��fD����rU4�m��g.�~�Q��g��ڰ��S��y���ϱ��|O���*Jw�)��Y��=R������B��+�n��NG	�L,�N�C9*�¢�"�,�>E���,�PK����Iihs[g��DW��ԅ1Qr��[��l_ ��b�FP&p�]f�"v!�`�(i3�5c�;�K ���l�;���EWrZ鎬����6�"����6ӹ%�ֱ�q��,��ur#��IH��*��B��<.+6J!N}�m��{�@��֯g�!�`�(i3Y%T��BP	�I]����2N��n��t�J�Yy�z�4�`�v"�,�>E����cfo�7>�����ǚr��yݶ�`�6#U����I��N}�m��{�������Q8p�=��[�зq8�Ј��{�W�%̷��q� �#�� �\�7>�����ǚr��y�7�cDtϫ���Uh1��:5A��p��èV����S`t�L?t����}>�O���(<�H�8�H�RtV�^�]�B#	�ƍ2���l�3���Z[�{�]��~9��c�	?�N����u?�:�H��$}�����U��E1tSjv�C���q(��v����om�K�w�H�<��wbk�$����$��-�	ڜ M�ݚ�Н����W��Ȑ�U���e��ݚ�Н��]��/ݐ=k_0�b�Y�{'%suE9�+����|��p�G	kp^y�,ԍQXF�S8�#�F�t��j��Ͳw���T!�`�(i3=aUh���P�|���9��V�9T�8o��7�Co7�wk��'���Xw
�T�r�5�ݑ���&�d>&S�XQ�?8B�����>a!~�)�=5U�i�J�8�7���}Dq�f��q�	��c0c �)��T�?�)�i�wbk�$����$���]�!������G��'T���+�#�C����N�DNl�q�#�-S8�#�F�t��j��Ug��d�M�}��,�)��w�19�"�����~7�X��u]yDy���W&�KKA�t�Hh�<LXn�tץ���:Z{G�i�e�n�^���Q�Y�<���%��ci���{2�wbk�$����$���]�!������G��+�t2������g��)�`�>a!~�)�=5U�i�J�8�7���}Dq�f��q�	��c�G�C�*۞���Yk��T�8o��7�Co7�wk��'���Xw
�T�r�5�ݑ���&�d�+��\���J��8��LS8�#�F�t��j��Ͳw���T!�`�(i3=aUh���`����	���SENan&���ߊ�ֲ���ܜ?n昼�2#:�^�V]��}>�C�;�����:=�� л���'��
���i�������l���=�64�+�E��&"�D'wg�������������G�R�u��r��!�`�(i3~�`cC�4��q�O�"pU
�T�r�5�!�`�(i3套�qD0��֋��V̷_��yC��S8�>c��6/�M��f�򃳿K��	�1��� ����P�7� �:5A��p�Ra])n#��'�ә�I,�D�y:��}���)��U�UH�RtV�^�y��j��k
�X�nZ�"��/B)�g��2���}Dq�f�<�6�Q=�G�)�<`�4];ˍH�r�W!k#��S8�>|��̂�!�`�(i3:�HCaIMl*h~U�?uӿ��hgo�I=���O�rs�i���(|�%%9��K�ł��
�T�r�5�
�:qEp<�@b`��%R�W"���z�X@*[�]�̵�7�!~u��r��!�`�(i3~�`cC�4��L?��.��nB_��j0!�`�(i3i`YS���2l�]<���������?�dh?v�!�`�(i35�����}YE+8�D��\���d��Q^�MY:�.ow�}l���Yk��!�`�(i3}A�4�/n�W�%cWʔ8k��.ͥ�H�RtV�^!�`�(i3w�����A��ߎ�x��y�g�5��zƍ2���l�!�`�(i3�����!�`�(i3�wӨj]h�O�M:R	�W׸���=C'�^�����ݚ�Н�
�:qEp�;�P�t�5!�`�(i3���W0�]��e|)0����n�=�Ra])n#���r�����'ѧ�Z,α�)IL��	�t�jGru
L�H��ɒ%Y$�~"Zr����fh����爮��J���ݚ�Н�$f��_Ub�F�S�1 ����W0�]��x@��m�ڨ�hծHN��R��bP�63Z�t�����
�:qEpbSo�3=�8���[{/;�;�P�t�5�x��8<��H8{�Fz�:pF��w��&���{[�����n/��dc�@c�����hfR��}��'{w#/ B��?	y�Lu��j��7�wtMM����+&�fg1c�:�(hS>�jV[$�)�vx4��<��^n�g.�5����L6�>P�2-i_m�;Y'�V1@�`�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�@hz�Rp�