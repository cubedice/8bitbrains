��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR�� (� ��"fف�����*z�w4G� ������[���a�8%`��4�s�6�XAoeu��a@����þ�V�\O����L�N��<G� �mD�?ea�8�����B}rs4������I���0�N<��;��� B]�pE���	x]̃Dj#^Da����M�$����o��I�绯�t�z����)�,�˛D��w���旴4w�1����h���������$[G��m$�;�`��v��p�㈍x���t�켻�S���c,31�-elwB(�93;2���Zߧl4���0�?�1~�x�c�>j����d��S�W�>��Q�d����t�mR��:�����-��3���7�Jk�b#Ӡe��?�F��&��q�©��7��#!l'���h�W�ӝ:X�{!�'�]��;�I�Qg�@zh�S҆�|n���,�l#�8�'�?�Tזi�!J�Й�m��8��r���t��U+�v��d���	u\��a(�m�Q� Q١Ӿ�$r�O��C��0��D�[T�Q~���c�K�$)���T�u���;���CXx��}�/mrH>pRݴ�c"�hf�7�o���R���=�K��%����\�4�sc�[�.���M��RwM���	ɭ8���#8�d��~�MUs ��?�L(	���&�Ll�ݍb�e����K��U�d?p�._q�l�2����v�`��H6�[	�V�D��~���pKJ�)6�X�e��D��8wɦU��D��)�.I�z���{����V���	x]�m�Je{q�F���S�V��R��.' J���<��:�%�+M��m}o����0���A����&���-Jv��k�8���҆�|n���(^k{3�)��t�����E)ԋ�J�Й�m�g/\}�����"��yА���k�9�N��U�o>#j~�˿_��h���O�`D��#�Bk�v,�ı{y�
� �AH�)��H��'�Wا[~�l]ǜ��*E����O�F@�4%���D�Pfc����2P����/�"��< ���X�M+��tc��P9P��`�.�D���J7"�x�YW��t��⫓���RL�a)3���ʉ�N	:.���n��Ex�W��"E`�{E�7C��H��n���`����A�dN ��>P�2-i_P�v�p�t,b		�����I� �o-�'�u�[U���z{��{k�DI<�m�����R@Q�V	��0NImh`�x�n�����w߽��-k��CG�)��h���
���g����y�=B<�O}=��Ѹ�7J_�:��r�O��C��0��$�>��wޥ�{%�a:���L����u���;����ڕ]��u��El��0{*r���8|�Z� 6,�0�T�vL [�AB�u�w+2^ݲ5�M�S��,�m~�}��0w�\���J�����\�4�s��{��]Qǯ�����շ��p��y�6율��'�~�MUs ��4ONw��9ӓ�t��^6ʯ*�a�WU�8s�#U�DN�9��b�7e�}�cz�m�!=�y����h�}`29�$zFs߬�����\K9�W��u���;����\_�MX�9�I�[��On�AN�.5f$��F�Ŋ�����}�K{ɈC`N�z����le�kI��Ř�^~tҦ,��_!���5�NnZsA���r�O��C��0���;f��jc#?���/� ��6�M�Q�8O �L#��&}Xa���qd��.�wjX5D	1�% �DZ�k�8���҆�|n����6f�@bU%x�eƐmt��߸I�0y����F@�4%��R�^�������o&��u��Uy��������RL�a)�ϕF���9c�J�M=���@"�X���-0�\8�:r&@$Y�q`�_����"��N�/��H.���{���}����X"��=��5�SK���Br�O��C��0��^������mߍu�M9F�*AJU��qχ�V���7C��H�j�?`%T=1�)�f�0��H��k3��Ԩr5@��_k���f0� �B͛	�m�O�����<�LZf4Q�����RL�a)	�n-�~Fc�J�M=�OSGM��n�ޘ���8�:r&@.ѿ)y�&���#����\S�W��`����I?�:���L�V$�"��D���i����	x]�fX�eϝ(˽0�9�(����-�[�D7n=�>��������V���8e3Z}�ax�� 5�k�8���҆�|n��T�{ ��ʥ�xw{���Fe����J�Й�m��/K5r�����}����Q������k�8���҆�|n���h��C dw�J�}d�j7n��h9L�W#�O�F@�4%��9��noM�6]3��|(*y�[oԓ�ҥ{E�?��RL�a)ѻtUWR����H7���[�(e��T~��)���7C��HʃE��z�ҷ�?�If㚍�4���zm�!=�y����h�}Y��݅ 0�)���K��Mx����o?�M��;]\V�A}��}���V���8e3Z}�ax�� 5�k�8���҆�|n���u� �(��)|#���{�`飨CJ�Й�m��C��ߊk'�4+.���`uI�[l٧cJ�^j�u��w)�S��X3���7��Mv�9:�A+�4ik"(�m"u4s8�:r&@�l�@��V1x�,�[ì���Tl��!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�
+&�s�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l����2�C�b��}Y���%�5�1�:�Ω�`<4}��)�Y¹w�yB-j&?��2�C�b��}�{b�2"���Bpш�#w��q�©���B���������'Sea�8���`<4}��(����5��4�l���+�Uz�QL<(�P[H�������'Sea�8���`<4}��(����5�2���[@%����nEAJ_�'��P9��6�g�m��+5z�P�_XV�>!�/�7��u���nEAJ_�'��P9�tw:g?�y��h�I����uk1i�f1?���b1�F��,��n�2��C�`Q���Ӿ���	���q��q�©��7��#!l'���h�W�ӝ:X�{!�'��M:��;6aJVlO/+�f�;�}�(�����_ q1j�iϳ��溂�U~܎VV����M��҇+:|8X����\�v�����Z���2��̪U��֜��3JHn��z�_c)���8�+�p}>&�&i���u*K6HT�����N��3w:��ݪ���`�����"IÙ=�H�ς.fOoI�J��#Kl�Y�7#�xI��Ok��@zL͊�q��UG�s�����M����A�m�(�� nU�IÙ=�HF���m¡��7=���bڕI��.E�b9����4�6�t�܀�(nԐJ*�Rs�08�b(���b9���P9b���a��cn��;���N�H}ة2�IÙ=�H%v@����fh�5,Wlr�r%)cA��u*K6HT�����N��2�F�P��U��+�Xa�H(�˕��u*K6HT�����N��2�F�P��U��+�XhU��`��&�b9����4�6�t�w�n����|��T�5�d�,W�� nU�IÙ=�H��'�PD����
q<O�n����9��#�B�sYC��\�v��_�R�G/K��(�������i{±�sR�{F;�f��X��Ye�?���j�g��$P�M	�D�$��띂ii�4];ˍH��T�K"
���d�8���obzĀY�ɡH�� �YߥթD�[*s��l=�L؅��FJ���/�`�����Y���÷uS�I0���ԏ�.fOe	m���h���b9���^F�Ј��m�K��� Z$���.>m�,kM:�yzL͊�q���\��;�,EfVNN��1��ݥ�U� ���_�ĕ|G���iyV�[g��� ��"��1��ݥ�U� ���_�ĕ|G���
�gγʝ�r6�>��/Z$�~�|Y�؅��FJ��� c�2��`���r'����<�=D��rMÏA�����i�؅��FJ���j`t���}Eo^������m؅��FJ���������ɰ�͝�e>����C8����̇i�d�?��E����F��j��\w��0]Y��
�iC"�,�>E����-��%Mό���.��6[��u�V�<�nbBIc��Et��q���U��^L��6�}�%b�CGފ����]�!��	Ǹ�y85����!��K|�d�MHOm�<G2s�%�8���/�l|�*"k���(ӈ���m�r����h��eZ�����E��@IE�U��>��l%i�-i��H�p�E����F7G#+��\w��0][�л���7"�,�>E����-��%M�rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0/v�K7%'c��Et�p�VU��Jm�QA�Q* q�\E��0</���/�u��(�
t��Y�{'%s:3���5C�ݪ���CyW�f�tR�wX��hs�����n��0�5	x��(�
t��Y�{'%s�h�v���&���$S�ݪ���CyW�f�t<|����faՊJ�e:[e��mea�8�����B}rs4������I���0�������Ls�F�%ܪ���PL~΄gO�3f��*����"�Q:�{�1��q�©��7��#!l'���h�W�ӝ:X�{!�'�W|�.Ҩ�$ BŊ���4��t���@H�o
��?�4b�$z@Q�:�ұ"��Q��4�2b6�e}�5����`K'�g.J/-ԋ6��v��o2�r��%��h,?�3�P��Z�N>�4�
����),��9��"!<<��u�	�sv�貛	#�蠿����66�v��G���V>�R<�2N��n���?���^��b9����{oS��n4s1�h�9�*�?�';:ZËF�3$����Vܙ��kE�{�N���0u�\k|aT��3G���"��y�S�yH��"J�A��S+�:G�W]�dט�w������Gl�N~)�jA( ����_�h3��{I��Z��H1c�f���2�خa�>����n8���ٳ��溂�ZI8'��@I��'��q�2�_:��p\I��� ±�sR�{F3�_� ��0���c�Br��VYW\_�B&��p���*��[w�'n�^0o�VU&ZM��9��"!<sB� 3�o`��K Yr��VYW\-@��F~*7���&�_0M�/�s���'n�^0o�'vX[��M�l��S�J*�Rs�08�b(��+�w]�B׿�ġ��,=�?���j��?� Zh�R?�R��ng.�~R���R	2͇��v�+ʢG&q^�`
�c��><�$�X~��\��|�^��
�>IÙ=�Hss2����`�|��K�z�H�MPq6.?�)���؀qjZ�`�|��K�z��|����=%+]Bo�A;h�F��O�i���AԢ�a\�D�����R�`�|��K�z���k��$a(􆿳��?ƾ�؀qjZ�`�|��K�z{�x���;�L���9�D_�3���U_�+X�܄�֝���b�Bϱ�����7���{r��I`1R�J�On`�(=�T�\ ��y�.�`L�
	�7F���I@1���t$I+�V�6IWJE�YY���F;�I�e�,��[�9q�Y�{'%s��.|Z���I7��-5��6��	���`y�����g�,P�n�Ͱ��Le�2l��4�y��ɦ�@^7&ģM�&yy��<:�W�_ĵn(���˧�0z�cUL3�X�j�>&�&i�"j���b7|#9����sC��I\�AkF˯�+)�Y�Q�d���'n�^0o<5�������Mj�(ȅ��Y^�@VJH/(f�|��*ܑe�W����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�����څ�ɡ��ls�u°������Г�����
iEE�Gr�ĵz��ݦ\�t!�ǿyXAm�Ln��S�W�כJϾ�ig()��ikp���H����Q#�?���;���Nå�a1����U��+�XhU��`��&m��1xс�ݦ\�t!�ǿyXAm��p�7 �s,�v����;^�6#9�H�MPq6.JHn��z���0+&�����|�F֣z>Q�Q�<%�a����D�K���g�,P�n�R<�����\���^�W+`�x�oP��@t�&�e�5
�`#_G�쵄����T�=�;^�6#9���k��$a(􆿳�f����DB�$��Xo��yذ��t�H�MPq6.JHn��z����#��F˯�+)���>�FFVx�%L�ib|� %�5����`K��M���-g?���ųJHn��z�F�x�aK�k����k!�\Z��K����C&��͞o�$C���8��'���ތ�1��\�vŁW�����+���LQ�$d`(���D7��%4������`-t"wdC��dט�w����j����r2��������������JHn��z�>�ack���A�;�֋`N(��/沄�J��CK��g�,P�nMN���OON�
_�n�@/%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7���i�_:�����k��$a(􆿳�f����DB�$��Xo����Ǳg�P�e�9��<���h��'n�^0o�'vX[���?� Zh�R6/��������рӚx��	��x���:%��Z���d���F}���3Yc�#�<�R�+}��hV�f����0+W���F�^�Y�7#�xI���|�r�HzL͊�q�������m	z1�Z���=�Ζ�,�Z{ �=�%��+y��yp�m~|�֙X�D��H�MPq6.JHn��z�%�,��CU���it	�TU����z~����.`Ϊ�/-T)x�?{���x.�Knq�]���7'����eR��x#2���p�����h��x�]�V���KD:�}��0nk��ކء�Ch�1Ǥ �)�?�0��Y��W���U�dP_\G�7^2$S�6���f�_)fxg��pH���0�Ҋ@)�t�d�f�rЄzɳ�B��,��C-2�^���ij�IROgn�t���c�&�<�o��H�,>��*�:��I�}L������@���t����N@<����fRD�}a�/^�yQA��D,��f�x��r
iEE�G�-��<s\�H��/Sg�w��'o��b9������|L�K�)x�?{���x.�Knq��H�����ġ��,�l�A���aZ��qA�E�nV�`=������!�`�(i3��Q]� _ό���.�}�
�?��]����w!�`�(i3!�`�(i37s�9���o��S8�)qcA�����M����A�m�([}�@��L}�
�?��e�S��@��Vd��· ���4�r�&Ɓ>i[�ͧ�?Y�f�kN�ı*�7`����\Z��K��4����/�����N���Q��B%Я��:��X�E����F�|��{�r�z��N��ξ���I��RhF���k��76����,D�+�8��io�iA'R�	:�@�F������L���a\Y���};l�-��;a���i3�|)sՀ]�N��&��v1a{J��bC�����Y��U�m?�o>����h�9��{lGD�V�B�x|qj0����N�}#�U��	�K�o�;*�}Ւ�~ܔp�l
d��U�9�r�<Uee�N�����H�OM��` R��B���gN�U�$etX��P��}�
�?��V5VM�dh-�kN�k�:A�	S�r��AR1<��J�@Ym��`�z��Y��),�B۸��L� s�j8����DzL�#�r��8��o[��ױ�*ܑe�W����n�4�`t��D����M����A�m�([}�@��L�@����gGKCYb,�q��iKXt(!K��tf��
_�n�@/%{�;����f�kN�ı/���^�"�k'	-����]�bgyvے�(�iF��׿]S��( �]�!��M8���	D%��_�ͅ������e����y
 <�1�����NĈ��r�]@P�B��X��8���/����,D�
�t�J8u���/	��:�a��Y�{'%s�[�&B�踫g(�r�N�ǁ�f�TIX����%V�����F˯�+)�"j���b7|#9���b!��u፤.��.f�Cz瀿3�7s�9���on�-�6��
�jW��D���M����A�m�(a?�X`.�-�ʙ@E>*;�¬pX��g��U-�e5/�=��kb!��u���j�4��(�[�*7s�9���o��S8�/ #O�)Ĉ��r�]@P�B��X��8���/����,D,Q�\C�8�Hj\��-��Ug��q���U��@����gG_$Mt�z�NG�և��f����Ր�z*���Be�2l��4��a��se�ξ���e�J�Pn\�pD��ZOUi3�|)sՀ2��2,��g�ܧ*y+k&v�IzZ鎬����
C��8q��f�kN�ı��U��+�Xa�H(�˕�&Ã�M�Ĉ��r�]@P�B��X��8���/�I����"�Oi9L�:�k]m��,�۞��	���/y��g�'b�t	�U���C��O]r�<Uee���R�}vJ^����`a��R<�����á�~O��L;Л��|#9���b!��u��Ɔ �����Vd��[�l\�`�|��K�z��@d��ץr�&U������G|M��i�ܰAb!��u��N�+k&v�IzZ鎬����
C��8q��f�kN�ı��U��+�Xa�H(�˕o�`�_f>&�&i�"j���b7|#9���b!��u��N�!�`�(i3��'�e��`�)�	�%{�;����f�kN�ı��U��+�Xa�H(�˕-+��B�Gh}Nw����=�����I|���bZ0!S�,��ш�A3�(N��㎏qló��@d����Q��O�بeD�I�Y�Q��*7b!��u፞�f
t斃����u_7s�9���on�-�6��
�jW��D���M���R'),��`��wu���뿼��8��''6���;8=�g��U-�e5/�=��kb!��u�]���!E/�x)�L�]�!��	Ǹ�y85�����5��d5�:�w�+���LQ���"X��[�d�a�4$�b!��u��D������������Y�{'%s���'����C�`�/�t��;mQ��8���/����,D��26N��-4e�[��]�!����w�Հ�	:ү0CAe[u�;0�7s�9���o�jƓ�[b!��u�L�������ғ�vq�\[$Q��
�̞��>���+���A���ۖ$����J�	�LÆ��E� )�&PW���[f|#9���b!��u��R=�"��ғ�vq�\[$Q��
�̞��>�˚? �	����`y����@����gGf���ѩj�7��'�b���b�Bϱ���w�K�1c+����Y~�y����u{ᵿ�����"X��[��Q[R�7ݓ��E�S���%��`��@�����0y�	 ���t��h�/a�'�̗�����C�M�����T�\ ��i3�|)sՀg�j*8a�.��� Ev�P"G�wk�١��	;q�ew�:��w�<om��F`���G���`y����@����gG��B��~7��'�b���b�Bϱ���w�K�b��2W hbvk~�#xTU]O�d��g��U-�ez�r�6��DP֞ M��V!�D�n`5�fK��0z�cULjaGkƊ~F˯�+)�"j���b7|#9���b!��u�+�uB;y�������Y�{'%s���'����C�`�/�t�KV*�3?�|��T�5�d�,WT	W $V��8���/����,DY�O�~H@1"�,�>E���]�!����w�Հ�[�=�5x��A~*aiqq��T���E@~����`y����@����gG��5�!�m��E����FZ鎬������_�,�;�7���c��չ�Ad��d�٣���N N�S�\�#$�ÙA�
M�<vW�n`5�fK�\w��0]b!��u�#� �,W�_�S�
ut�q���U��@����gG�0����Oid�w4ZxZ鎬������_�,��|[p2e�F;p�	�j}"K���rs�i����ej1W��Mw���1�Z���=�"j���b7���Øf}�
�?��I�_Pg<�l��姹�g�YӅ:��U,�(�)8���0y�	��sC宸I))����A�m�(/!���La|#9���b!��u�G9�:Q��Ĵ��ޯi�ʌ	���bSq��T�ٮ|�,
���]�x}NI0���ԏ�.fOe	��q��"o��Q[R�7�)�`E5�j�W��� D�cg�}��E�`JcUȵ�ixUS��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ��i3�|)sՀCeFJ5x�_�k]m���E��Y��(���G
\[$Q��
�̞��>��b��v݋N��������(($��R�wX��}�
�?�Q�>�H�(�{��U���!�`�(i3�U,�(�)8⋌�U2ރ�8���/����,D�Ĭ}��򛚆z�Ji�!�`�(i3y��Fp����f���,(���B����Ӝ$��BS�>�!/�_�n�To�[
MQ9�F�����#oM|#9���b!��u�[��m�U����#31�#��d_O�=�ͦ�١��	;qS�>�!/�_�n�To�[
MQ9�F��g��U-�e,%�0g���j�|�{'�v1a{J��7G��D@���B+AԢ�a\��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ��i3�|)sՀ*�şxˏ1��o\�B/�`�B7d���lJ��튝�b�Bϱ�����7���{r��'6���;8=�g��U-�e,%�0g���j�|�{'�v1a{J�j�f�At�a�W��f���,(���B����: ��ao.\C�kHgN�����`y����@����gG��l��`��Ĵ��ޯiڡ�F1�4W1�c$^f42�|�,
���]�x}NI0���ԏ�.fOe	��q��"o��Q[R�7�����bp�WdM4@��_�U*�D|[H�%"ȵ�ixUS��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ���s!�k�����k��#��
��\(^Fn�H�~M�"�,�>E���a�x���w�K��f�
l�w1�����\�H��/Sg�w��'o��W5OL���I/J}�
�?��֗�_{h�!�`�(i3!�`�(i3�k�XLF�<�rם4�S��ł�!r�1�Ѯ�a�}�
�?�K�\7}�W,��+G���tJ]J�a:��U,�(�)8g��dT�W/S��8(�E���Kt����ӯIJ ��`y���h}Nw��諚��y�[�l��姹�C�`N���Z.��0�W\[$Q��
�̞��>��b��v݋N������M}Ĭ���1����X�[��`y����@����gG��l��`��Ĵ��ޯi��ŁO��8�P��Ά���0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX��}�
�?�K�\7}�W, D�cg�}Ŭvc��W�ғ�vq���q�41&q^�`
�c��><�$�X~��\��o����׋��`y����@����gG��l��`��Ĵ��ޯi�d�A~y��Fp����L�de��-@��F~*7���&�_���/���l���F�8���/�I����"�Xt��R�F��6�ғ�vq�\[$Q��
�̞��>��3
�v�v-}�	mp�?IK��y�8���/����,D�KlAP}k�`�B7d��U,�(�)8�}�Y�ןw�8���/����,D�KlAP}kScmWP���U,�(�)8�K�o���,�z��f�|�?��t���2����.〧I����k]m�����i�#Ѻ\[$Q��
�̞��>��b��v݋N��������(($��R�wX��}�
�?����D)���Z� ��(HxZ��j�
�&�j��1�a-���7a
��r��L;Л�����Øf}�
�?��I�_Pg<�(y�.
جH?���)xZ��j�
�iB{�Z�_�1�����\�H��/Sg޶��j�}a�cfC?�Q䨈��Q[R�7�)�`E5�j�W���yͧT���E"����5�Wȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e,%�0g����]�gv���J�����/t4S��]���f���,(���B����: ��ao.\C�k�ף�D�~�z$��8���/����,D��ǉã1X�v1a{J����nFy� ����Uҫ��0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX��}�
�?��I�_Pg<���7�*w�^Ϗ�'�xZ��j�
�iB{�Z�_�1�����\�H��/Sg޶��j�}a�cfC?�Q䨈��Q[R�7�)�`E5�j�W����΂o����^�?�ȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e,%�0g����Ed��>�^�v1a{J�"����5�WúAV�!s���0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX��}�
�?����D)�ܮ�S�Gz�!�`�(i3xZ��j�
�&�j��1�a-���7a
��r����~v����"X��[��Q[R�7�
�CӞD��m�q�/��v1a{J��Z�n�f��AԢ�a\��F�dH�/�O��� ӫ/��m�A0`��A1Q"(L��8���/����,D,Q�\C�/�����	^%�R��tCtHC�'Ϯ|�,
���]�x}NI0���ԏ�.fOe	m���h��D�P�E6���2����.0��jOT��.m��TDZ��O$��lJ��튝�b�Bϱ�����7���{r��I`1R�J�On`�(=�T�\ ������q�f@��L���N�b�'Be��-���AԢ�a\蟖�S� ?�0��E|�,°������R�wX��}�
�?�N��	�Ȓme":l�n�U,�(�)8Q�y�� Y{q����'6���;8=�g��U-�ez�r�6JL���Z'#y�>�)L��H"҆>X�¨�Rk�6�3
�v�v-}�	mp`g�_��iB{�Z�_�1�����\�H��/Sg�w��'o�D�P�E6���2����.JL���Z'#y�>�)L�/|w~S."��*Ha���J*�Rs�0�ǳ7��y.�k�XLF�iB{�Z�_�1�����\�H��/Sg�w��'o�D�P�E6�ټ*w2�56�)�`E5;]MBg2Zr�G� YF��6�!�`�(i3!�`�(i3!�`�(i3�E����F�f���,(���B����: ��ao.\C�kHgN�����`y����@����gG�7�{�mo5i,�Ĕi��)��ۺ��fyd�F�O����!�`�(i3!�`�(i3O�=�ͦ�١��	;qS�>�!/�_�n�To�[
MQ9�F��g��U-�e,%�0g����]�gv���9$��i�Yi䚠疛!wFii�"�/̯��39�#c�ᜂl��=5;ى�,
_�|���0y�	��sC宸I))����A�m�(/!���La|#9���b!��u���a�vw����~m�(��k8!�`�(i3!�`�(i3!�`�(i3"�,�>E���a�x���w�K��r�]�4�P�l��=5;�<��|��k�8���/����,D��ǉã1X&U;��]�x�'��x!5�kz���[h�b��v݋N������\!�ZJ�k�XLF�iB{�Z�_�1�����\�H��/Sg�w��'o�D�P�E6���2����.JL���Z'���V��H?Ә�%"Q�ܦfM� �L�Y}śT�!�`�(i3!�`�(i3зq8�Ј\[$Q��
�̞��>��b��v݋N��������(($��R�wX��}�
�?�rS����u�}�Q���GM�о٫�]�r�Gפ ި�6v ӫ/��m�h��"��ȵ�ixUS��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ������q�f@�]�gv��JeYSWe^E1��b�����=�?I®|�,
���]�x}NI0���ԏ�.fOe	��q��"o��Q[R�7�)�`E5�j�W�����ד*(�E��W�u&�Pߺ0��A���ۖ�s;�Ê�\[$Q��
�̞��>��b��v݋N������M}Ĭ���1����X�[��`y����@����gGQ��6��'A�{�>�� ��
�m���+)x�?{��
0#`�1��ȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e,%�0g����]�gv���J�������ߧj@Q�_Y��t��3
�v�v-}�	mp�l��U�h�|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�|#9���b!��u�G9�:Q��F��P�?��4�+��_碍�(H0et�?����0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX��}�
�?�G��-�HG(�b�'Be����\)Pߺ0��A���ۖ�.Q�2�>�f���,(���B����: ��ao.\C�k�ף�D�~R��v	�R�wX�ո@����gGQ��6��'w/���h8%L�瞩w�jȐ���,��a�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ���sC���X!�`�(i3!�`�(i3�p}8�JL���Z'm&����T�ˣޫ�B��i��)��ۺ��fyd�(��|Q9XI�|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�*��/qRr!�`�(i3���aR�}�
�?��I�_Pg<˃�B�1Yw�Yi䚠疛!wFii�"�/̯��3�{s��ֹԚ���$\[$Q��
�̞��>��b��v݋N������M}Ĭ���1����X�[��`y����@����gG�6�
}St� ��
�Q�
w�8F��6�O�=�ͦ�١��	;qS�>�!/�_�n�To�[r��}k:�~�ȧq�6a(􆿳�����r9E!�`�(i3���aR�}�
�?�����4R�ت����¿'��x!5�kz���[h����XzR����(ZAB���0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�Г����ѼmJ�0�6�b!��u��!�jT7|�`\%��u7W�:����p�A[wN�hH����0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�Г�����!�`�(i3m�ڨ�hծ�)�`E5�R(R�X���Ǹ���m�(��k8һ��6��b��QM!Ϊu��U)�ȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e�,���6+��dט�w���[X-�BM�ܤm|��Z�j-J���\�v���eQ��`��ļަ��P�5��/dV�z~~�Y_"R�W�uw�2�w7u>(����r��o��])x�?{���x.�Knq���e�-yH����8�YM�S�I))����A�m�(�$��&w@}e��(I0���ԏ�.fOe	h~S�O��}�6[�O�?�n�� <!�HI9َ���vV6\PJ�x;����#��2歮/"Q�r0�Z���s<�>5������֐^�݉ ��|�`q�L��S�E!Sb��&'��G�,Bճ��s�l�En	ғ�#�O+�� �ד�]#����z�Ji�ғ�vq�\[$Q��
�̞��>��Z�<��H��h �=�����#oM|#9���b!��u�Y�)�}��EXs70��lJ��튝�b�Bϱ���w�K�	�<���BSG�p�P��<jV���\�H��/Sg�w��'o�6��T���7�8���/����,D�>: �.�� n2ϒ���=��pA( ����_�s�G�J�;�s��&<����A@��CazrZtc�!{p85��Ph���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�Q��VC��.��Ԟ-zq_��Wj�)I��-�q�1f]�r�r��J G3͐j8�&?-��{O��c_`J��Y��)�.����ktL�j
�"��d���!iS�4F{+�i7N�_�Ar��� �Q��ǺΕ�A�m�(���
�u�
_��s�֙7�}�!��]�0^ݵT";��|BP72���6�������c����c�QN�~lAW,u��#7���>�Y:�{;�s�c��K��Ƕ�W�}�o�Z���@	�<����$���D��8�tufJ*�Rs�08�b(����X�zgz�'�̗��������,Լ�Se���7�}�!��9�{�Jj3�a�5@�i��V,'9k�6!�`�(i3J�a$�Y �+�ϸ�i�	��+@�@�VҒmͦ���ҧ�GR�D^f�Nd+l�Yҽ֗�51����~��`Z�h�l�Rk�X�Q��ǺΕ�A�m�(慧��a���}Dq�f�����,�ǰTm�v��G�6��~p�=��$*Im���O?a.���J=R������~��_T���a�aq���)�F��Օ��qvdЧ^{�j�RtW���d���!i�wӨj]h���6�ü��k>B2�6�zX���+��T�����D3���������M!�`�(i3t�iZ]XF�hx��G��!�`�(i3��x��&^�B�wj$g�X;p`�ct�:��RE3z%�u�܆!�`�(i3�����ݱ������]�`�g()��ikp���H����>�#P�'�̗������צS0��ݚ�Н����8��T�h���}둮j\����C��rR#K�p�ݚ�Н��K�^��Q��G�S>\.�!::tm�0�i.�9!�`�(i3eX+��f J�"e~��O��!�i�3���j�\�"����ݚ�Н��� л�|�9I����o�u�/!�I=�+��2Y��kک�x����y���ݫ�ф���F�)!�`�(i3���ȍry��	�B�'��a�F�,�U6�Q�L��!�`�(i3��0�&�ͭ�U젩`#�4>?� �1!�`�(i3��"����M몴PBoT�ݚ�Н�?V��j�c�
���!8ϟ��7�4�Mzuf�?ǉ�=�2��}���zgm##��V5VM�d6��0]�1�v�9��s->m�9V��Vv��8>�=������iG��Ӆ�+��T�����D3���������M!�`�(i3t�iZ]XF�hx��G��!�`�(i3��x��&^�B�wj$g�X;p`�ct�:��RE3z%�u�܆!�`�(i3�����ݱ������]�`�g()��ikp���H����>�#P�'�̗������צS0��ݚ�Н����8��T�h���}둮j\����C��rR#K�p�ݚ�Н��K�^��Q��G�S>\.�!::tm�0�i.�9!�`�(i3eX+��f J�"e~��O��!�i�3���j�\�"����ݚ�Н��� л�|�9I����o�u�/!�I=�+��2Y��kک�x����y���ݫ�ф���F�)!�`�(i3���ȍry��	�B�'��a�F�,�U6�Q�L��!�`�(i3��0�&�ͭ�U젩`#�4>?� �1!�`�(i3��"����M몴PBoT�ݚ�Н�?V��j�c�
���!8ϟ��7�4:i�P.j*�7`����\Z��K��l�W@i�!�`�(i3{k�h�+d�/Y�Z-u�}#�U�����Y)N���������$��@�n���I��)���W�w��fDV�o����!ݲ��_)�d�h���{w���z��(����5���ռ�j�ŋ������Dua�\�:��)giR�7h�,b0V�u�Q�ݚ�Н��w,�����<v���G�=���Q{�1�a-���7a
��r�,���9^-�W���`moF˯�+)Ƌ��_��F˯�+)��&�C�/L/���?T�x~1�@��@�Ce�<�˹�40<~�>b�eIG�5�}�]���p.0��I�!z���.M�ݚ�Н��dv��oTN֢&@��&Zt%��m&<	.������Z鎬�������(���ڔ6�.���Vd��S��g�lE!�`�(i3%$1�q���0��"��S8�TkF����v1a{J���
]$�P�v	��Y?V��j�c��99�)b�+5�4��c�YC��?�!�`�(i33�kM�}��s.�֡m�\�&e���
�s��wӨj]h�0)xU����V5VM�dj��;q+#Cxz!B�`
 ֢����oC������U{a��f�?ǉ�=�_F�k-�H��bf�?ǉ�=��|��p8=�[Ǵ��p���@Z���%>�rG�<�]�Ե�8h�7w^D��/��iG��Ӆ�+��T����oGo�Z�K����ހ d���l�6>8G�%?gV��U�x�l��1:�N�*�x��'T���+�htO!��nT�Ā���-@��F~*7���&�_j;��q,!�`�(i3w¹��<d�Ji�];���w¹��<d�,��L��!�`�(i3n�NQa"_�?���C[u��oŹQ!�`�(i3EfVNN{s�ܱ?'�EfVNN�����1I^�e����kn4@Q�/�!�`�(i3�EhP�Q�ug�%Y��̗0z�cULj� 1��k]m����� ���*�7`����\Z��K���Pxە���!�`�(i3�%=��Lg�%Y��̗0z�cULj� 1��k]m����{"gY*�7`����\Z��K���Pxە����ݚ�Н�[�л���7��{��W�����A@�Q��ǺΕ�A�m�(�]�	��f�?ǉ�=q�\E��0���N��t�3����_�Ξ)�N�ǁ�f�TpD��ZOU	XT�1�wӨj]h�0)xU����V5VM�d|�v�W��I4��欱���j����,X�|H*�ݚ�Н��9+��������i��W��¹���I��RhF�� ��*�C�ժ*)xJe��hy��)]W��7#OOJd֯�y��j��k����U{8�C,0�?���!�`�(i3E�l�����5Ƈ���	I��)���W�w��fD2�e��P���x�NS$x���z*�7`����\Z��K��itXgWZ�G�+5�4��c �&A�5I��RhF��F4#_�h�L�R��k9V��	��y:�^c��D`���J�.�$`b��8�>r&�N������8�C&y8_��s�֙4�(�Ҁч�+5�4��c!�
�!��V5VM�d��0�8k���;_��8W�w��fD���4�-lT��{B�z��z6Y�m@�<����I�?g�f��Qө}�_g�?�H���w�1#fr�L�t�iZ]XF�hx��G��Zt%��m&<9U:����VK�5��&q^�`
�c��><�$�X~��\���.x9�S{���2��̪U��֜��3�F�7��Y�
�cc�V�x��7��0�趦����'���o���a5��I�~�џ0I� X�1���g���}| ��+qѭ�+g[�|�\m�� �8B�@`6Y�{'%s���F����:�#�.��N�x%؋��LrÁ���G���%=��Lg�%Y��̗0z�cULj� 1��k]m��d�r����ArCcGXO�P�v	��Y���S�|J�s.�֡m��z���_ΩI4��欱���j����u���tt��2��}��6d��H�_�ϟ��7�4y��4��U�*�7`����\Z��K���9�u���=?V��j�c5;���0�+5�4��c�H�v�m��Y��)h��{���3��� �Rmu(�������e�-3�i��7u�`��Y��)h��{���Y���EP��_F�k-�H��bf�?ǉ�=��:��"7i�m�T�੉��%>�rG�<�]�Ե�
'��u���*ь��MᖡtWKj���lJ����I�?g�f��Qө}�_g�?�H���w�1#fr�L�t�iZ]XF�hx��G��Zt%��m&<9U:����VK�5��&q^�`
�c��><�$�X~��\���.x9�S{���2��̪U��֜��3�F�7��Y�
�cc�V�x��7��0�趦����'���o���a5��I�~�џ0I� X�1���g���}| ��+qѭ�+g[�|�\m�� �8B�@`6Y�{'%s���F����:�#�.��N�x%�UZ���s����G���%=��Lg�%Y��̗0z�cULj� 1��k]m��d�r����:�繇q�P�v	��Y���S�|J�s.�֡m��z���_ΩI4��欱���j���֬���[pq�\E��0���N��t�3����_�Ξ)�N�ǁ�f�TIX����B7Ԅ���ra5�k�K�s.�֡mh�l�Rk�X�Q��ǺΕ�A�m�(D}����4�/�"����=�m<��_2jV�T��I4��欱���j���֬���[p�_F�k-�H��bf�?ǉ�=��:��"7i�m�T�੉��%>�rG�<�]�Ե�L�J~�H�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��"Jc�l�!H��R��M��gq� �ɰ����Mp��Q�V��&��C5YD�H*�r�wl�({�x���	R�N~)�jm�w���i���Z��FkH�������h	�(����5���&<˴m�TJ	V�+�PM�^-q�x�l��1:�N�*�x���N�4���f�����Q�_f�Nd+l�Yҽ֗�?Mة�1Zn����������\����>'���������6%�a�<çI� yMŃ�,��) �?��7��qp�ToJ�Eyz?]4�f�?ǉ�=�m�n���֣��n��ݜt���,\ͨ܉p����O,8�ݚ�Н�bs��2[������	�;�ݚ�Н�0q���Q�L��
�:qEp3?���*�YmC,igu?V��j�c<�s����	��7��u���/	�C\�2x���?V��j�c�?�#B,��	��7���=��ծ�C\�2x���?V��j�cZ)[���F	��7��z_nÑ2h����>PҝbYގEV�kn��KG*���D5�|أͽgF"?�Q��ǺΕ�A�m�(It8Z�QC;��|B
y�3~;�>ۀ��t�~x��	��#�c�'����������Vo[���˚����Z��L�{	�����p�� �&SfzF�.z9��+5�4��c~�t;\p�I�{�P������ j��U�`��d�Ϲ�r��`Z��\�&e��\'�s!���I��RhF��L>�/�G��g��b�w�R���ykb>���pۀ��t�~x�_��.���n�8�Z�Ѽ���9$��H��u�d�ۋI7��-5r�p =(��8�B���ow_;O
�J��:�����7��|qAܡKy����nFW�JyS�.��.f���T��M5�*5o]E�HN��R��?�d���&��_$U����-�߃�}����,�ǰ����
k�=�w�x�Șoj&P*\�m�ڨ�hծ����,�ǰ>�l�s�wE�=p���u%�RAo�����igu���_r�e~5�O�%E#P���S����i7N�_�z*K��I4��欱���j����Eo(d�J��:�����7��|qA�&+��`��51�X�c�rs�i�@24b��H�[���wk����E�E�L�t��n�"+n��,r�I7��-5�������K�i���r������,������u��XJ6dq�e$ct�:��RE8���168Ow�R���yv4�����=��ܦ���u6j�"Hs�����{F��w��s2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>�����J�uT��&�Zf`��"����h��^�`�����t�T��?E-h��`f���sd�G}%����3f�'w�4�5wFlE� ��'ž1�|�'����u��r����@�z]���ߋ3]2dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&rG��Hb� h�ҩ��T�T�y����S_��̷_��yC��S8�����ZK����E~��G���۵z �+5�4��c�H�v�m��Y��)h��{���=e�0S��D�I7��-5�������:5A��p���F��O�}�	76�&�� Ӗ�t$�)�vxn]ϲ8����Q嵉�edy"���h�v6�z'kKǹ|���|u��R� l���E[J��:����b!��u���j�4�<�..�4�Ὗ�i�#Ѻ'���Xw�j�7�����$�/���$ڿ��Fյ[+8��a8r>yP��b�G�lnO���Tq��A��sp!!v*!�����m���pQw�t���o�eW-���C#/<���q��c��qVw���lŀ�<J�Rz��j�4�¹��� Y[� ߨ�1�� ���E�N���n�WP���9�űW��Cr���v�_���!I���?ML�˔?F��v_}�S�Z��tb{�H�C�_�Z��{a�g�Gc^���Hxq"���w[	zF�F�=��� *	�Qu�c5rQ^5�y���3Ve�
w+B$4IA��w����=R��B�"}��o�u�/��Bqz��9��daA��Cm��mἨdh���b�S]���o"83��Je��v»M�{�|Lɣ���d��TD��5��b�Bϱ�H�^B�3�A�'�.����PԹ���!�`�(i3!�`�(i3!�`�(i3`
 ֢���XƤ5_��,\��ݝۺ������M���X�^��D����jVѭ@!�`�(i3!�`�(i3!�`�(i3��7I���&�<���8}
��5-���:)�
�9��W�&]�6�o8:4�I���c�90B3v�A��{y����i�q,?5q��7���9��j�4�<�..�4���|#HK��A(�c���_G��Hb� h�ҩ��T�T�y�8�Hj\���i�{ypP ��j�4�<�..�4��G��}X��?��t�-=���]	"e��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r��Dw\�����b�S]���o"83�� P�jc�8�Hj\���M7#� �6���n6��dh_��tC}ߟ�r�Q��b��Bgk"������m�q�/���e���W�.�]ؔVG��"X��[��Q[R�7���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}ī��K��M��y��{�"���b��Bgj��i�s���j�4�<�..�4��C&��b�:)�
�9LeQp�K֣����[$R�i�Yl-H�1O�N�
w5���iѕ:�,�����4�G-rx��� 0v��W5�WIi{4D+G��-�HG($R�i�Yl-ҡ"#�k�1���~!�`�(i3!�`�(i3;�x'_|~�뽢�7;6ik!�S���{ �4"-��/��,�Q��M���I�m�J���z>9�R��d���!i��$o����8��lq%`,9�H�W@�kr� U����n�j�Q��tf�á?�d���&��ݚ�Н��:�,��f!��������raǹ}���,*r��@�VҒmͅ.�g3Zꢯ�wv��QX�mR�HN��R��?�d���&�(���o�����-�w�R���y��}���mD�W�G�ZL�]�2�.�|���"FS�_
���.{Π��yGb�:"�G�}��d���!i�T�T�y�8�Hj\��/�Y��x�!�`�(i3J�a$�Y )P<�ܓ�Y��9Ӌ�L`���(�oh�5,Wl�/�O'�=�s~`WGW}ߟ�r�Q\ b�{�$�P����9�oh� qs��l��v�`,9�H�W��`�z���n�j�Q��tf�á?�d���&�t�{#	�x�}�������IЫ�Is�8�w\�PPO�s"�6
��E�i�m}66j�"Hs�^��rWI
"d\>�7��U���V��	��yIV�q���t��^�T����Y����S2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�I���Y/�/�hǙ cX�d��?6��H��X�����k楊HaU$kX�M�ŗ\�'	�?��[n8�A�A���p������'HY-��Yk"1/|sL'���oֲ󄰊�������M�����%kR��������֢&@��&���o)�]r k�|6�8NU�:|������k!�\Z��K��f�?ǉ�= k��%�ෑ=���4��#o�;-;*�7����E���=�<���� zL���s�`���A.o�G�m�?��x�Mu�W���`moF˯�+)�H�f�M�&�����ϲ���6%�aj:�Mpp�}�(�-l̜	H��d˹�40<~I�~�џ0I� X�1��kޮ��g��� ��"aJ �!,|�8��5ǛHO��E��������~G����EX��dC$,\ͨ܉p����O,8�ݚ�Н�K�\7}�W,:S�.?<N��	�Ȓ�@{2귑�7��m�K�!�`�(i3+�uB;y�e����'�N��(���K�!�`�(i3I��
�[��b=��y��j��k����U{8�C,0�?��ʉ��%>�rG�<�]�Ե���5R��T��t]�<Lz+M�ᴰ`�V��rU�w�⽒��8�>r&���R�}vJ^�k��76�;��|B
y�3~;�>�������\t��r��X9���R<�����á�~O��#t:0���nS�3�ǻ��d���!iЈH�����b�'Be����s:��Ϲ�r������D�v1a{J���V!��N�$r�t�}iV��	��y�� �P�qN+M�ᴰ`��_��.���9�Z�y�6nZ:ӄ��8����"O��o���ia������v�h�g��U-�e a⣃_B7�}�!��b8IU_h��Rhy�������D����u_�*5o]E�HN��R��?�d���&��|��Li�8j�H�p�.�g3ZE��g�Hb�t]�<Lz+M�ᴰ`�dТ���S֜���,�ǰ�+9\���������������>�ܫWEFΑǜh����X "
z��_r�e~5�O�%E#P���=J����uS�#̮y�3���;_��8W�w��fD�1�C�#�] �y�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�"��3E9�H�i�e�}�������B�@o��[ea�8���	�~����a��+��#fr�L�t�iZ]XF�hx��G�����=�-�o&l������g����=�tt"���O�����J��a�U"�������o��\�l�Ϧ���I�:뼥<7.��H�ʱˡFZd6�o�·���~X�~���$^!!�`�(i3uwТ�
2������}�k�+9=����Kp&�@���k��-��w¹��<d���	fd,���9^-��כ��p܏�<
DN��X;p`�Vx�%L3z%�u�܆��O���R�^Ƒ��!�`�(i3*bL�(R��u��n�k|p��z~���8��'@���k�� tZ�u���ߘ�)�Ij;��q,��
4#!���ڃ�"�!�`�(i3�������t���ck��,�:�N�*�x��0�&�ͭ-��i�m�T�੝�hy��Q�#<4^�>N0Θ��;b�-�2�>c��?Ӈa�/!O�f�?ǉ�=�<��>��%@��4��).i���SRX$��V����覭L��G�dE�h�����?�O̀���vj��$��覭L�q�\E��0	ozqPx�6_s/��g������n3�x�h�k�t]�<Lz�l#�V��H��<�C�Ar��� f�Nd+l��p��;z�_��s�֙R���Bk�d*e��\@8GS��`n������ct�:��RE�QS����>�wo��Z��Ac<�p{�5�O�%E#P�P����9��g�ܧ*y*J�X�$����aV}�������,���1����,H/������,�ǰ�������'����2�,bxqX��g�9��,Y�����9C�������u8q��ǵc��5�%]����8�B���ow_;O
�J��:���闺����ő��"�\�!�{~����DKY�����|f���+X�E�k?�i2�.[W�w��fD�g�9��,Y��(c$�,w�R���y���,!��HC�d��g���'N3 �zY]�埅�t�į��>�n��-�U4��\w��˪?�-�l~�U�n��(���_��s�֙R���Bk�dNmyM<�G�ۺ�Ub�!�V��u��i�_:�����k��$�8�B���ow_;O
�J��:�����A��AC�m]���z2�nFW�JyS��f
t斃����u_�*5o]E�HN��R��?�d���&�c�����|�� 7�G�Yw�R���y���,!��HC�d��g�[��f��*�)|/P2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>���yn�4^4 ��#�$G�l����M���R'),��`ތ@�'��|0;��|B�v��䣞�a���~�(����5���&<˴m���q~�i��+��YR�7h�,b0V�u�Q�ݚ�Н�}�\�����nW����p���,��2��������")d���ݚ�Н�w¹��<d���<
DN��-a6@v�+U����z~���MK�LS�_�p���it	�TU����z~���3O�)���_�\G��4�	B45j;��q,G����?���_�\G�k�y'��a�o�� ������it	�T!b%�ZV�p����nZ���t��˳3[�u8�̇i�d�?��X;p`�l.�	�C˟B�'��a��7��r�=H��bf�?ǉ�=�|�)՜�4�X;p`�YmC,igu?V��j�c>ݣK�6<oC7z����f
t斃����u_f�?ǉ�=�� ߌ���X;p`�]���!E�0䇙[�v`ͤΟ�}a�~~��}H_��i�;��%YM�	�v�3�2������"�*o�yG�f>x�:	Yk�2�4.��̈́��3R&�5�V��X9���i�_:�����k��$�8�B���ow_;O
��ۈ`4�`1�����j��G�m���*J�X�$��¯ԙEI�s+��6�.|th1�$�g�O�M�,*	V��	��y�� �P�qN2�W1S�]�tH���]*?�d���&�zY]�埅�,Ǥ���(��/z*q+6j�"Hs��zX�k�wE�=p���y2Z��Zk���T�}ɻ���}J�|���|����wC�5'�O��d���!i!q��V��������pĀc��ŏG�m�����C*�	�V��	��y�bB�.���O�4��ϐ!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��_~�TP�[!�� Q�N6l��F��#cj1�g���(����5�Z��f��Ո��D��2E#fr�L�t�iZ]XF�hx��G��n����������������i�����d]���GF��a�1�Z���=�,���9^-���M���R��ӟ-��<P��C�Y~�y����6d�dG�7:������a�^��D��j��&��8!�w� wk���,���9^-���0)]��w�b^X�P�9���TE��a��'�-�1H�3}�?�_�������� "5�]֭�h��Oo��0��7t�%�Z?��<�ry^�h�'f R�X;p`�(������\�LtF�&8�,�#N�)L�*�_�I<�N��KPkqy�{"�i:�gR(]ͅ�y�����5�.?V��j�cB�Y���c
=�2����޴�ik]�)�^�\�� ߌ��-���h��=;��bC����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�P{���b�������IQ�%�+2�}R���
�f�<�vd�̪ǪzAV:Ń�}M:y8s�1E���7������I�R�ω�9A[1Z��`��!��>�� �ڬ������F ���Ru���$-�Hq)��p�����R�Zm?�QgS�
 ��baC`֓�5��/`�#E������.#f{}#k���P��#��s�'	�?��[�-���^��Up�OSg.V����7X���8C��D9�C�W6r���["�=�bB�#fr�L��ϸ��#|S������3[�u8��� ��w��]n���І��%n3������k�+9=���(��U��֜��3�AQ�0G�C�`�/�t��ߖ Y��U���gFck
�������}g�2Y��kک����n|�p[Y���"����)�-}�|ݔ�3�z���.Mp����nZ���t��˳3[�u8��M�g����H��bf�?ǉ�=̇i�d�?�4�0 L?�p���@Z�6[��u�9k�\,���K+!q���!�`�(i3扈�[-�c]^�mOeTky��2��}���zgm##�+��%�k<�^�V��	��y�3�&A��SwE�=p��-:�N�Ò�}kutC������i{��*ȑs;��|B�Տ� �*��q�)�`C�G����]'\gWg��	�Z�kfc?�#	*]]�(&�L�xjzӝ���I(͂��-�����2��}��cVe�U2�<��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�G`B� �'����u��r���2��}��cVe�U2�< 'J��@�D`ks�F⽉��%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}���Q���!���ūaT��3G?�d���&�s͟;)f���KXL6�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9Y���&���'܍|Cy���QJ�wk����\����|ݔ�3�(n�'�(�S��)��R�^Ƒ��;��|BEΟ��
�U�a�(��^GѬ�_���t�T��?E-h��`f���sC>��ӚH�RtV�^�'ž1�|�'����u��r��q�\E��04>^!b!4b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3��Nh�=f[���������<�.�����8��GM��-����!�`�(i3�v�Wס���G�K$x/��&���PC-��i0Q�͹�Ɩ,�b�R؅�!�`�(i3q�\E��0����G�t���m�� �ݪ���CyW�f�tR�wX��!�`�(i3��Ě�����}Dq�f��3��C���H�� �YߥթD�[*�Bi�v�V���;AD�e�{�W!�`�(i32+5�"�����-P��F����~�;2V-W��	c@�^ k�R�e�0���m�e#e>�=�^݊<���He�ylB��-t���m�� �ݪ�򈟕��+�v�7��]�ݚ�Н�3��0����g����F����~�;2V-W��	c@�^ k�R�e�0���m�e#e>�=�^݊����xQ�e�ylB��-t���m�� �ݪ�򈟕��+�v��t���?�� h�ҩ�!�`�(i3�lTN��I���q�}���{BO���5�%]���a(􆿳����^��!�`�(i3��jVѭ@!�`�(i3u?�:�H�jsrCm�k�J��6�d�t��w��X�'����u��r��!�`�(i3q�\E��0��@Z���rs�i�}�O��LTSG��ʎ�=U9��R�^Ƒ�Ӆ��I�ѪtR�^Ƒ�ӆ�v�9��!�`�(i3�����!�`�(i3�wӨj]h�(%����Z鎬�������(���/%Z�ڄ^1��#ƌ/B�ݪ��2�r5�����jV�{+�fbmDF�!�`�(i3���%>�rGO�D mWN!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ o�n�J-�ƪe�0c�)�Ul����,�ǰ	r�R��Z����i�|7��_	�s�t�{���6������]'m���G�K$xE�p4rqG7]u��
�3�R�^Ƒ��;��|BEΟ��
�U�a�(��$��,Ix�6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3e�v��ҵl�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r��pT/�GS��%�����d��-��![L��^C�+a��o���H�RtV�^q�\E��0��@Z���rs�i�@24b��H�[���wkL�1p/-��G�<6�U����z~)���	6�
�:qEp�;�P�t�5fĉ>99��A0ok�׹�3��܌o��oŵE=��X�z��V��	��y�߬9�6ש�ڔ*��T�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc
M����n��i���~+�lX҉ޖ�˞,cƶ��^�}���8�\�(fw���I��RhF��0��N�F�6��9I�u��'����(fw���I��RhF���,�=R�/��Se����-���^��U���P[�񁫴}2��uR�9$��i����t�T��?E-h��`f���sC>��Ӛ��S�J\7!c�2���j"�²O�y���0ܔ��'ž1�|�'����u��r��N��r8!�k]m��Z�����hh��,��Oˊ��C����t�ǊS�>�!/�_�n�To�[
MQ9�F�1�m+�D8�̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*�Va�ir���M��2"���&�^��v�8:?�'��ᦾ�;���8���U�._�nQ�rV��q�t7�v�]��1���U�._�h�5,Wlr�r%)cA�r�(�%�pH�RtV�^N��r8!�k]m��Z�����h���G��S:t�L)��k]m���E��Y�^�Mi~_�T���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�������c����g��U�S��q�}��il���iA'R�	z�#,gB��Pߺ0��A���ۖ�)�-�W���a�x�G9�:Q��Ĵ��ޯi���l`Zd�g()��ikp���H�����[��l_G9�:Q����v�z`���ө%�Sg()��ikp���H���׾ŞWsuz��"]c�#y�>�)L����0ˮR�m ޶&�hbvk~�#x��#�H��+���42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!H�x�7X�J�����_�U*Cw�Hm���9��N	{8G9�:Q��Ĵ��ޯi�I#�(���)x�?{���x.�Knq^nї�Y�_�n�To�[
MQ9�F�����
��\�H��/Sg�w��'o�v��؄aX��I�_Pg<�l��姹���Mt��a�x�]c
j���l��姹�ȃT����A���ۖ��S�<Ԣ������f�l��=5;֡Q��Ⱥ���>��� ӫ/��m�D�K��D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�C�7ª6��J�����_�U*Cw�Hm��G9�:Q��Ĵ��ޯiڼ�ze��>տ�:
hbvk~�#x+[.Sk�NA�I�_Pg<�%��g:�����<�ׅ��A5W��v�8:Tr�E	�[��J�����_�U*��ө%�Sg()��ikp���H���^?������X��O���r����!�`�(i3!�`�(i3!�`�(i3�I�_Pg<�%��g:�����<�ׅ��A5W��v�8:C��4�I[��I))����A�m�(�-4�{>��G9�:Q����v�z`�Cw�Hm��G9�:Q����v�z`���ө%�Sg()��ikp���H���GM��QО#y�>�)L�/|w~S."��*Ha���J*�Rs�0��|�_�Y�j�W��� D�cg�}��m���+)x�?{���<m�N=-�w���+ާ�����ݚ�Н�!�`�(i3!�`�(i3 #��zG���J����k̇���APߺ0��A���ۖ�èr�L��b��v݋N�����&r�"A��A���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9g�O��B~��0Ր�5Ҹ�u�����φ��<�6�@a� ��fFMqlgd�G}%����3fUi���Z�͗�M9f��;�jmT�#bs��2[�a��o���H�RtV�^�}��il��o\�B/�k9a�S6��_
�u �V.��$��l��=5;r�$�(��{�R���/�O��� ӫ/��m8D����#U��,H/���k��^�1��dc�@c�����h��-����;�jmT�#�,l����?0G.{T�2��^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���F�H۷`"��]ap��e��>��Օ��qvdЧ^{�j4�����ݚ�Н�޼QE1��v1a{J�)�H�b�b�Bϱ�G9�:Q����v�z`���+_AdV
�:qEp�;�P�t�5fĉ>99��A0ok�׹��*P�{���"��\��}g��V�;ܬo>v<~<�=a��0� ޼QE1������m�(��k8!�`�(i3!�`�(i3!�`�(i3!�`�(i3+�F�$-�S:t�L)��k]m��l��e b6vJ�pZ� 4�F�Α��Dr�2�N��r8!�E��Y��Q�
w�8D�t�%o�V���-$�!�`�(i3!�`�(i3q����`U�0�V;�M�J�����_�U*���$����;-�]�pR�$5iL�Pf8e���N��r8!�E��Y��Q�
w�8D�t�%o�V�g�yl��6T�T�D��ao.\C�k����S�{؁C�*&#�4?�o�5�h�B�c\��L̎C��fx'v�ao.\C�k*h�!<^Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������Mڷ���o\�B/�i
�i�w�Qטg�u2�Tt$Ó6N��o\�B/7� :(c�Wh<�!C���>��� ӫ/��mo��7�^�1n��y��a3G7```+��)_�32�K�y؄@�!�`�(i3!�`�(i3����&��+�%�t�*#y�>�)L��H"҆>X������*fW� �/88n
I��jÇ+�_�n�To�[
MQ9�F��,bxqX�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcU�۩}�w��k]m��
ae���K�9�*��� c(H޵D7W�:���iޚuq6p��j����Q�9�|`ЉɁmwlc(H޵D7W�:���k!��,�<��y�@�v,����.�u-�w���+kGA��ݼ��r����!�`�(i3�o�5��!<��y�@�vFn�H�~M������f�l��=5;O�R'o��!�`�(i3sU�@{Q�p��j����Q�9�|`ЉɁmwlc(H޵D7W�:���k!��,�<��y�@�v,����.�u-�w���+�\#���Ƹ���r����!�`�(i3���>�t�mo5i,�Ĕi��)��ۺ��fyd�,m �\��\�H��/Sg�w��'o�'uFէ���p��j�����8"c�։Ɂmwl�E��Y��Q�
w�8D�t�%o�V\�Z�0��9$��i�Yi䚠疛!wFii���_�?2��HL�U���W�H�2^�/3!�`�(i3�0�9&،�d�G`5[��{#Ÿ�&Sq�a"��ř�!�`�(i3!�`�(i3!�`�(i3�����wP?��i/R�c��;=~. .����mo5i,�Ĕi��)��ۺ��fyd뉯ӌ$/k�&U;��]�x�'��x!5�kz���[h�x�1W0�-��4��Ɂmwl�E��Y��Q�
w�8D�t�%o�V�g�yl��6T�T�D��ao.\C�kT���/T$�&U;��]�x�'��x!5�kz���[hin5�҇�?�b��v݋N�����U-�pë��";Yy\'{w#/ B!�`�(i3޼QE1�&U;��]�x�'��x!5�kz���[hin5�҇�?�b��v݋N������G������p8�Iט��ō�Zm\�l��ì�A؁C�*&#�4?�o�5�h�B�]�{����d�G`5[��{#Ÿ�&Sq�aM^�ؾiZ-�w���+�gVdxQ,��a�vw����~m�(��k8w��?L�@���wp>�\�H��/Sg��'|F��d�G`5[��{#Ÿ�&Sq�a���y*/@(�_��%$>_�n�To�[���&YH��-��k���H�2^�/3!�`�(i33��0��e��0�U+�qbp@��C�7ª6�9$��i�Yi䚠�5���u�L�!�`�(i3!�`�(i3!�`�(i3��c���鿉�X+�kQ��v1a{J�i�\��ou#���3qV�[�U�b(l�rD��ЀUg]�6��;b؁C�*&#�4?�o�5�h�B� ި�6v ӫ/��m�h��"��^����'5��9$��i�Yi䚠�@CF���(�b��v݋N�����&r�"A��ArS����u�}�Q���GM�о٫�S��wE\�!�`�(i3!�`�(i3�I����~u͘6��q���j�W���]�B� ��8@��1�*)�2�"��wb���E�¸>`!�9wY����<��y�@�v�&Sq�aj(��;����_��%$>_�n�To�[�pI�
KrS����u�}�Q���GM�о٫���^O�K����fx'v�ao.\C�k*h�!<^Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������Mڷ��iA'R�	��}E-��$@PJ+5*�轓�A1�J�����_�U*����e��ھC��'#���fx'v�ao.\C�k C�Mh�n �O`�Ag��ۭXX�|ʡi�����Fz�!�`�(i3!�`�(i3����&��+�%�t�*#y�>�)L��Bѭ�pR�$5iL�$�F�V��&|���BY��l��=5; �e� ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���Mڷ��iA'R�	��}E-��${`�9$��i�Yi䚠��&���)"r�DyA�S⏸[����LG��&��a�vw����~m�(��k8���wp>�\�H��/Sg��'|F��d�G`5[��{#Ÿ�&Sq�a�_��%$>_�n�To�[���&YH�HL�U���W�H�2^�/3!�`�(i3�0�9&،�d�G`5[��{#Ÿ�&Sq�a�_��%$>_�n�To�[��H	X�ʁ���Mյ��#�@����ۭXX���E��O��d�G`5[��{#Ÿ�&Sq�a�_��%$>_�n�To�[B���v��؁C�*&#�4?�o�5�h�B� ި�6v ӫ/��m����	���γ~<�����6Bj�!�`�(i39<��`f;]MBg2Zr�G� Y� {l��	z�9^Ȑ�I))����A�m�(�W[����p8�Iט��ō�Zm\�l��ì�A���V��H?Ә�%"Q�ܦfM� �'9�5���c(H޵D7W�:����p�A�ԍ'8�����";Yy\'{w#/ B!�`�(i3޼QE1������m�(��k8һ��6�!�`�(i3!�`�(i3!�`�(i3�����9�Xy+�Mk��趵��1�F���������m�(��k8һ��6�D��)��	u�}�Q���GM�о٫��s�~�L�1{&��� )S���z;]MBg2Zr�G� Y� {l��	�g�yl��6T�T�D��ao.\C�kT���/T$ǩ����m�(��k8һ��6ݕ��wp>�\�H��/Sg�u-Y2�G�1{&��� ���xl�ݚ�Н�!�`�(i3�V3���L�瞩w�j���@ΙN�[���-ل9�#c�ᜂl��=5;J5�#Z�"r�DyA�S⏸[��t��7�M~�V3���L�瞩w�j���@ΙN���HPԎ��V��H?Ә�%"Q�ܦfM� ��x�1W0�-��4��Ɂmwlc(H޵D7W�:����p�A�z;#o"�I0���ԏ�ʖ�:���V3���L�瞩w�j���@ΙN�[���-ل9�#c�ᜂl��=5;� Ek�0��������mo��jVѭ@!�`�(i3��dN���ub�z'hۉ)��_�2��|2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!��7&���Y'=�t%�!�XH��Oi�HU5��)4�3Yb�J+c%F���_�z<���L1v�}7>�W��	2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��:�dy�v1a{J����%]+a���G����E������7D!��l��姹�xAQ�Y;x����̜�I0���ԏ�.fOe	���X�a1p��j����Q�9�|`Ю�K49AԢ�a\�[�U�b(lƿWdM4@��z(��xo}E�٦���sC宸I))����A�m�(�QNȮ���k/��m#ׇӭ��!�`�(i3!�`�(i3h큈��{��UJ����"]c�#y�>�)L��H"҆>X�(JdT�ݙڈ�KK?B�&�_j����)Ł�I��jÇ+�_�n�To�[
MQ9�F��(��&��[��m�U����#34�?��˧+P"G�wk�[�S��]c
j���l��姹�I�oൠ��ڈ�KK?B�&�_j�In)0LH�* �b�p�Ĵ��ޯi�-Qq��Pn���G��(��{�O�iA'R�	��}E-�c��n�#&|���BY��l��=5;\�Z���O`�Ag��ۭXX�|ʡi������ڈ�KK?Ba���$_Ĵ��ޯiڡ�F1�4WM7�FM\�1�����\�H��/Sg�w��'oª���#oMA�H4$B����>��� ӫ/��mt�����W�br�*7�iA'R�	��}E-��0��ٟ�͘6��q���j�W����+G��ܻ�ߣA����Dr�2��c���ğ�%��g:���
A�%�q����	�����͘6��q���j�W���]�B� ��8@��1�*)�2�"��wb����,]�������ڈ�KK?BD�1N��λ�g��ZR�,��9 �ubK���E�g��ZR����z�Ji��1ʟÛm�w��ГQ�H���&�b �hvT�+]�x}NI0���ԏ�.fOe	-=3�$��ϐa�x�����on�b�Bϱ�m�(��k8����~�䱢�z
A��Φ�gz(AٸI))����A�m�(JX��!�.�`;���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcq�(Ul��?U�D�K�X�K{�(��	}�@�r�<Uee�N�����b��[cS;��|B�V���p�e�S��@��Vd�uҹW3�"b!�`�(i3!�`�(i3�s���6�v1a{J�o1J����٣�}��iA'R�	�z�?��D@N�ǁ�f�TpD��ZOU���Gx5��WdM4@��_�U*�>=:9_�aV��	��y���x.0��X��FO��(���*�`�
��pF泥���k2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ᾣ4��L}c��ko#k��^)�Qטg�u2�Tt$Ó6N��o\�B/�&���+��h<�!C���>��� ӫ/��m�D�K��D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�C�7ª6�JeYSWe^E1��b���S�C���0�V;�M�J����'",��X��a�x��"�%�U_k���$,@����:_��k]m��Cw�Hm���V3����C��z��&���)"r�DyA�c(H޵D�ҏ@n�k!��,�Sc��h� ����r-�w���+kGA��ݼ��r����!�`�(i3!�`�(i3�V3����C��z�ob.�Y�2W�b��v݋N�����&r�"A��A���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9g�O��B~�z5�0P�ġ��x���u�Y�KG�ξ���I��RhF��F4#_�h���Se���7�}�!���e�S��@��Vd�Y���DO�!�`�(i3!�`�(i3a�u��e�MN*�������*y}e���:�#�|$.@L�`f�Nd+l�Yҽ֗�51����~�gKh���V�H�M�I��)���W�w��fDl2����}*�NRcnvyw�R���yW�R�w���L�>5�C��Ҁ"���`Vk�d��f�Nd+l�Yҽ֗�X�e��n�ސ����U��)���Y;e�iK!���d.���+�^n=\f�5>�HҰ±�͹�uR�:l��xjzӝ���I(͂��-����.[�Kδ9����˦G�K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н��I��� g~��q6g�yF}���V6l;�<��'�̗����Ep� �����4br���^��D�Ϛ�-����!�`�(i3�P�궊�2�����8!��?V�ы�(�)x�?{���x.�Knq'ێ����� h�ҩ���6��5=��)Q��h�xF墣c#���K!�`�(i3�����!�`�(i3Zi=���lr�{��|e��0�U+�qbp@�!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ�d�n�ͻ���~͏닓.�`�3���M��,�IX0F�MV�ҁGG%4vkz����`���φ��<�6�닓.�`�3�P���F\xjzӝ���I(͂��-��������FYs%?es� e��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����M?��y�!�`�(i3<�g��H��&�2���)x�?{���x.�Knq��5+*��d�@���G�X���.��ġ��,��5+*��4br���qP�V>t'�̗����S]�_�_��u��r��`
 ֢���֦�n��{_8�Y��=�}�Vݨ��}Dq�f������!�`�(i3s�3r<��AgC�&��������5�,D|r9�g()��ikp���H����m-F���T�YN
��)e���T���b�Bϱ�h�5,Wlr�r%)cA�5QN���d>�c�n�P3�K��b� h�ҩ���6��ZRR����Mn__���q�Ӯ�!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�MI8�ѐv2Q{VcҟA��0Ր�5��v/�(%줄$�HY�����A$�P������5d��n4s1�U��B��-�*P�{��Ɖ�<�(]|kY-�xjzӝ���I(͂��-����N��r8!S⏸[�nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r��u?�:�H���^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���Fie6ӭkk�v�]��1���U�._�h�5,Wlr�r%)cA/�r�]/2�ݚ�Н�޼QE1����"���dN�<@Iv��nt=:��:5A��p��w�w:�!�`�(i3^()��>�����U�._�h�5,Wlr�r%)cA�r�(�%�pH�RtV�^M�yx�,�G��i/R�c�${`G7```+��T�TN��!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�M��uR3��%<�X1H�w���ސ����U��)���Y;e�iK!���d.���+�^n=\f�5>���u����uR�:l��xjzӝ���I(͂��-������T��xW����˦G����P�|T�T�����U(���B����Ӝ$��BS�>�!/�_�n�To�[
MQ9�F���v�9������g�Z��3��a���!@�f")u��r��܌;���'����u��r��u?�:�H���^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���Fie6ӭkk�v�]��1���U�._�h�5,Wlr�r%)cA/�r�]/2�ݚ�Н����cJ�C����o�W�F}���V6w��EO"�̞��>�_9�R�5;�/�O��� ӫ/��m�QP�*Hd��:5A��p��w�w:�!�`�(i3"G���RG7```+�ֶ������YN
��)e�W�J��H����8�O�5���1tSjv�!�`�(i3pR�$5iL̻��Fd]�ob.�Y�2W��C�Y�\�fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹��Li�AE��� �Rɴ��S��)�5���sO�v(�y��U��)���Y;e�iK!���d.���+�^n=\f�5>��UE�'���(0̈��N����"sS<�0�zG�������&G #��zG���J�����/t4�q���o�F}���V6� ��=y�̞��>��b��v݋N������M}Ĭ�����Gf�߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����?0G.{T�2��^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���F�H۷`"��]ap��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3G9�:Q����Z$�x$�֯� W(���27:։�X+�kQ��v1a{J����nFy� �ֿ�JO���%>�rGO�D mWN��Ě���aT��3G�IX0F�MG9�:Q����D����1����ciAG9�:Q���O7�4[i�$R�nS�]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7!c�2���j"�²O�i.����bs��2[�a��o���H�RtV�^G9�:Q��Y����(��U� �,\���͔5��:m�\�H��/Sg޶��"���̺`����1�����\�H��/Sg޶��j�}a�cfn��ٙ��Z*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81-���7,D|r9�g()��ikp���H����m-F���T�T�n��a��#�GWW�<om���m-F���T�YN
��)e�W�J��H����8�O�5���1tSjv� #��zG���J����0;�������G1=��͘6��q���j�W����΂o����^�?��:5A��p���F��O�}�	76�&�� Ӗ�t$�)�vxģ��_�ڑ8�`Lv�RU��P��i�u�}��il��J��O�����!�o��_�Rv�䩲$��8��I�:Fa�7���W"�P�K�0_f��3%�~eG���A(�c���_G��Hb� h�ҩ��I�_Pg<�(y�.
جHR��o�W�,\���͔5��:m�\�H��/Sg޶���W�Z[��MQ�'���1�����\�H��/Sg޶��j�}a�cfn��ٙ��Z*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81-���7,D|r9�g()��ikp���H����m-F���T�T�n��a��#�GWW�<om���m-F���T�YN
��)e�W�J��H����8�O�5���1tSjv� #��zG���J�������ߧj@Q�����&��"]c�#y�>�)L�^b٫
z�(;-ob���;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��I�_Pg<��4���Lo�h:E�,�do2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��PdG9�:Q����Z$�x�vG��*Ha���J*�Rs�0�ǳ7��y.��c���鿉�X+�kQ��v1a{J����nFy� =�r��J*�Rs�08�b(��g]�6��;b#y�>�)L�b�@_	���UH���4տ�:
hbvk~�#xo�������Qטg�u2]c
j�����7�*w#;���W��m ޶&�hbvk~�#x��#�H�޼QE1��v1a{J�Bz��s�V��m���+)x�?{��
0#`�1��׾ŞWsuz��"]c�#y�>�)L�^b٫
z�s�ť���)x�?{���x.�Knqo���n[�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE���Q��I�_Pg<�4���TS3���/k��1x�a��2e�>���x��j�W�����ד*(�os}�&à��b��v݋N������M}Ĭ���.�f���I�J*�Rs�08�b(�����̜�I0���ԏ�.fOe	m���h��v��؄aX��I�_Pg<���7�*w��D��q��S�C���+�%�t�*#y�>�)L�b�@_	��)�p��ZI0���ԏ�.fOe	m���h���s��訌��v�8:������fI��jÇ+�_�n�To�[r��}k:�%��H�7���|ss�j�W���yͧT���E"����5�W9a�Fc��Ǔ��K��v1a{J��¸�k�L�����f�l��=5;R�ˊ	18��X��g()��ikp���H�����V1G�׊�b��v݋N������M}Ĭ���E�����{��D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�C�7ª6��J�����/t4"����5�W�����G�v1a{J����nFy� �_Y��t��3
�v�v-}�	mpÊ�����j�W�����ד*(�E��W�u&�Pߺ0��A���ۖ禡�Q���#y�>�)L�����/s=s��4�+��_��A5W��v�8:'w/�'��γ~<����jVѭ@!�`�(i3!�`�(i3!�`�(i3 #��zG���J�����/t4��UH���4տ�:
hbvk~�#x����I0���ԏ�.fOe	m���h��g]�6��;b#y�>�)L�b�@_	�"����5�W�����G�v1a{J���Ꭓ�[���ө%�Sg()��ikp���H���GM��QО#y�>�)L�b�@_	���UH���4տ�:
hbvk~�#xa��H9��k]m����\�6��_Y��t��3
�v�v-}�	mp�dA�M}.F!��D�����k$ !�`�(i3!�`�(i3!�`�(i3�}��il��A�{�>�� ��
�m���+)x�?{��
0#`�1�������f�l��=5;R�ˊ	18��[	�"~�}��il��Rm�㭼�S}�S��� �~�^#y�>�)L�^b٫
zܫ5u�q��	�����aq��uG�բnG9�:Q��F��P�?��4�+��_��A5W��v�8:Tr�E	�[��J�������ߧj@Q�_Y��t��3
�v�v-}�	mp�dA�M}.F!��D�����k$ !�`�(i3!�`�(i3!�`�(i3�}��il��Rm�㭼�A�!�[��5�*Ha���J*�Rs�0K=X���d���fx'v�ao.\C�k�ף�D�~����Jϑ��+���42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�؈G�j��m&����T��Ŗծ��7W�:��e���b�!�`�(i3!�`�(i3!�`�(i3q����`U�0�V;�M�J����0;����0
"8�'o�*)�2�"��wb���E�¸>`!�}��il��G����1�E�AvY�5�h�B��A�	���\!�`�(i3!�`�(i3�I����~u͘6��q���j�W�����ד*(��j�Y|��a�x����r͖���"��Id�fPa[��I�_Pg<˃�B�1Yw�Yi䚠疛!wFii�"�/̯��3�{s��ֹ圂�Zd��(̚N�:R�j�W���<�'��V�I�'��x!5�kz���[h�\�n��I0���ԏ�.fOe	m���h���,bxqX�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ᾣ4��L[��m�U/|w~S."��i�*O����Qטg�u2R� [�'a,�v1a{J���Ꭓ�[��[�V�+�6f6,�#�I))����A�m�(};l�-����!cI͸I))����A�m�(};l�-��?�%�'^ȴp��j����Q�9�|`��Y�m�k?j!�`�(i3!�`�(i3!�`�(i3|0u�ښF���A�k]m��5L5@�m��B��رzh4�+7{�R����� ӫ/��m�A0`��A�"��(ޅ���>��� ӫ/��m�A0`��A���/j)	 ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���Mڷ���o\�B/N�.�L�0Ϩ �~�^m&����T��Ŗծ��7W�:���iޚuq6p��j����Q�9�|`ЉɁmwl�F��M:J�5���d��!�1G9�:Q��HN�YH8x|?Ә�%"Q�t�ч�����mo��jVѭ@!�`�(i3�� 3�m&����T��Ŗծ��7W�:���rL��7�_�n�To�[r��}k:�>�hy�!�`�(i3�ݓ�W���"r�DyA�S⏸[����LG��&G9�:Q��HN�YH8x|?Ә�%"Q��(�K��F��M:J�5��,����.�u-�w���+�\#���Ƹ���r����!�`�(i3�VR��)Đ�G����1�E�AvY�5�h�B�͞_'Bi��fx'v�ao.\C�k�ף�D�~�ڭRyԍ���#�@����ۭXX�WŚl��E�j�W���<�'��V�I�'��x!5�kz���[h'9�5���)�5���sO���%�$�m�(��k8w��?L�@^?���W��j�[O����k$ !�`�(i3�}��il��G����1�E�AvY�5�h�B��A�	���\!�`�(i3(*�O�q�@��i)&
�k�����oT`kz��{V�-_8���G�7W�:��G�z㤧{�>
�eEQZ�G����1�E�AvY�5�h�B�ˊ��6Ԩ{�1{&��� )S���z�j�W���<�'��V�I�'��x!5�kz���[hin5�҇�?����XzR��M��e��)�5���sO���%�$�m�(��k8w��?L�@�b��QM!i�9�s��^?���W��j�[O����k$ !�`�(i3�}��il��G����1�E�AvY�5�h�B�$5z&�D���ME�R�, &ấ<b�(*�O�q�@��i)&
�k�����oT`kz��{V�-_8���G�7W�:��G�z㤧{�>
�eEQZ�G����1�E�AvY�5�h�B�ˊ��6Ԩ{�1{&��� )S���z�j�W���<�'��V�I�'��x!5�kz���[hin5�҇�?����XzR��M��e��)�5���sO���%�$�m�(��k8w��?L�@�b��QM!i�9�s��^?����8������k$ !�`�(i3�~�7p����nt=:�+�_0c �I	�����g[�s6{޴�i��)���1�#��d_!�`�(i3!�`�(i3����;q�a�x�G9�:Q��Y���g��{�6G�a�x����r͖�k���$,�C�7ª6�L_v,<=��}�I����&Sq�aQ�y�QF��fK�Ěk.!�`�(i3^����'5�L_v,<=��}�I���Fn�H�~M�y�)w��W�l��=5;R�ˊ	18��[	�"~�qi4�747B��[�<?Ә�%"Q�ܦfM� �L�Y}śT�!�`�(i3!�`�(i3+�F�$-�S:t�L)��k]m����DބiMb�R�f��a��;���=����qFz�}o*o޼QE1�Bz��s�V�r�G� Y� {l��	�g�yl��6�����������iv�!�jT7|�`\%��u7W�:����p�Ǎ�͚�3�_�n�To�[r��}k:�b�	.�� ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>ht)PjL��k]m���E��Y�"����5�W9a�Fc���F���A�k]m����\�6����~�	hnp�����b��v݋N������M}Ĭ�����V1G�׊�b��v݋N������M}Ĭ���N��E�Q�>�H�(�#ve
��e����R,�!�`�(i3!�`�(i3!�`�(i3��+�t2�a1�����G9�:Q��F��P�?�?$٭n�rD��ЀU�r`�JtоI0���ԏ�.fOe	m���h�����̜�I0���ԏ�.fOe	m���h��֕ߝԀ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��4?ڇ���WdM4@��_�U*�^�?�9�*��� ��\�6��#P��Ѐ�N�w�qX�f��EJ,�G7```+�
�HYF�@�����4R�ت����¿'��x!5�kz���[h����XzRL��MWX��\�6��#P��Ѐ�5�h�B��ME�R�, ��Ѻ��	�1{&��� ���xl�ݚ�Н�!�`�(i3I	�����g[�s6{޴�i��)���!D������eW�d/=me�%b\%sU�@{Q�p��j����Q�9�|`ЉɁmwl��\�6��#P��Ѐ�5�h�B��ME�R�, m��
~�B�H[W2q�[�Kx�ʁQ7W�:���|���~�Fȯ+3�YE\����oW�l0����'{w#/ B!�`�(i3l�[K��K8��DބiML�瞩w�j���@ΙN�z�}��b��v݋N������M}Ĭ���N��E�p8�Iט��ō�Zm\�l��ì�A�����5qo��o�����&Sq�ae:rmv�H�!�jT7|�`\%��u7W�:����p�A�ԍ'8�����";Yy\'{w#/ B!�`�(i3޼QE1�Bz��s�V�r�G� Y� {l��	���-$�!�`�(i3!�`�(i3�����9�Xy+�Mk��趵��1�F����Bz��s�V�r�G� Y� {l��	\�Z�0��)��%��+b�O~1��GM�о٫��s�~�L�1{&��� )S���z�R(R�X���Ǹ���m�(��k8һ��6��b��QM!Ϊu��U)�Fx�Ǻ^U�:Q��z�˔ �y=k�2�u���e�՝*U��eW�d/=F�[$��<���H1���~!�`�(i3N��r8!��DބiML�瞩w�j���@ΙN�[���-ل�{s��ֹ�Em��r�~�����wP?��i/R�c��;=~.T"O5�`�7B��[�<?Ә�%"Q�ܦfM� �'9�5�����DބiML�瞩w�j���@ΙNVB=�4�S�-��k��[�����������5qo��o�����&Sq�aj(��;���Q�y�QF�靰v j}�!�jT7|�`\%��u7W�:����p�AE2p��Fȯ+3�YE\����oW�l0����'{w#/ B!�`�(i3i��r�+�<�W�.�P�@���?���"'�nH/#���J�ďx'��I�`�
��pFC�R��<:�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcU�H8����2[QvA��֣T�5��$@PJ+5*�轓�A1�J�������ߧj@Q�h�%��?Q_�n�To�[r��}k:1x����̓@?5���嚚3�%�I))����A�m�(};l�-������l�Y;2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��0<�$#y�>�)L�^b٫
zܫ5u�q��ҏ@n�$@PJ+5S:t�L)��k]m����DބiM��pqo�}�;-�]�̓@?5��l�ҵ�_�k]m���^�?�9�*��� �k]m����DބiM�YG5`FFB5=��)Q�n��y��a3�J�������ߧj@Q�_Y��t����M���X]c
j���(y�.
جH��O��U
h�07�;|''ZT��*�/4{+�x<�;���jVѭ@!�`�(i3!�`�(i3M�yx�,�G#y�>�)L�^b٫
zܫ5u�q��ҏ@n�rL��7�_�n�To�[r��}k:�b�	.��Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �b��D�씴SZ���U��)���Y;e�iK!���d.���+�^n=\f�5>�Ml`�`\Ձ���� \���F�`yx�>�+X�M?��y�Dw\����.m��K�+���w�c�c������_
�u϶=f�'�1�����\�H��/Sg޶��j�}a�cf�Lͷw���]�x}NI0���ԏ�.fOe	m���h���%@{Ex���k��^�1��dc�@c�����h��-�����s�Yls��8��GMm�HxX����U�._�3
�v�v-}�	mp
���U{���8^��hJL��;���N�4��N	�7q������O�޳!?�R��nścp�B��-/a8V�Ո���m�q�/��v1a{J��a`p�W�8��b�Bϱ���j�4��k]m����,^�V�:5A��p���F��O�}�	76�&�� Ӗ�t$�)�vxMl`�`\[�H�l�b��D�/�����	^%�R���m���+)x�?{��
0#`�1��9a�Fc�����^dE��C�x!�H��SW]#��5�m ޶&�hbvk~�#x��#�H����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcx�dŕ�n��.m��K�+���w�32��B��Qטg�u2c&��n��C�x!�H����'^_J���"~6���aq������n}L�I))����A�m�(};l�-����!cI͸I))����A�m�(};l�-������l�Y;2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���j�4��k]m����,^�VC&��b��Ɔ ���Ve��˅���ө%�Sg()��ikp���H���>��B�K�.m��K�+���w�?�H$~��	�����aq��[��n;�D/�����	^%�R���m���+)x�?{���<m�N=���fT��F*�L��!�`�(i3!�`�(i3!�`�(i3;�x'_|~� �S���}�cЉ�M�+!�j�8�3
�v�v-}�	mpl�!����_�n�To�[r��}k:�b�	.��=��5a�y�iA'R�	:�@�F���,�
�CA_�G��-�HG(�b�'BelĈ�\פ��
y���)_�32����r����!�`�(i3!�`�(i3!�`�(i3�G%�MP3ö�3���:b׻���3�v1a{J��bC�����'�NKc�F�*3��ö�3������7�V�k]m��d�r����dQ"��؆��)x���l��姹�-��#��e�S��@��Vd�2 ٭H�So	.���T`A�WdM4@��_�U*:J����#SX>tG�zi�X�+2�ꎷĬj����M��v�}졞���$U������h�̯#DC���C��Wo9����4~��E���ZaL݊���2�"�G�p�Pڹ��/^�w?�d���&���5�G
m�D ML:�N�2	�����8�5�IX0F�MV�ҁGG`5:�����+�^n=\f�5>����5��M������S������"sS<�0�zG�������&G��6���2[QvA�΁�a�n���I����~uK7͍��|��W&":�ݚ�Н����D)�ܮ�S�Gz�J�a$�Y dN�<@Iv��nt=:��:5A��p[�t��#��l��姹�g�YӅ:�E�g�������(ӈ���m�r����١w��zj�v1a{J�&��	�>�n��>�my$�N��o�/���;�/��@���WdM4@�k̇���A�C��|uK7͍��|��W&":�ݚ�Н�K�\7}�W,��+G�����̑:�dN�<@Iv��nt=:��:5A��p�T�T�y�/������Z� ��(HE�g�������(ӈ���m�r����ЈH�����b�'Be΁�a�n��n��>�my$�N��o�/���;��6�����
y��!�`�(i3�I����~uK7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv���6���2[QvA�΁�a�n���I����~uAԢ�a\蟴���P`��ɠD(c!)��w�K��r�]�4�P�l��=5;���o�1g��U-�e1�S�������6���2[QvA�LO�>��
�I����~uAԢ�a\蟴���P`��ʱ�O��W���]�x}NI0���ԏ�.fOe	m���h������#oM��:<��j!�`�(i3�⒍~����v�z`�!�`�(i3���G��(��{�O��o\�B/����~�(���B����: ��ao.\C�kf��_@Z��T�\ �͆�v�9��</Sn���k]m��Z�����he�an�P�ݝ�b�Bϱ�[��m�U�H"҆>Xĭ�����̞��>��b��v݋N���������L+-�8���/��:5A��p١w��zj�v1a{J��9H�P�.�}6�/S� ����,��WdM4@�k̇���AG��&'��̞��>��b��v݋N������M}Ĭ���F`���G��k/��m#��}Dq�f����Mڷ��iA'R�	z�#,gB�������&���e�S�[�k]m���E��Y��%�i����w�K��r�]�4�P�l��=5;R�ˊ	18?.���|�T�\ �͆�v�9��Dw\����.m��TDZ��O$mQ��RA��m�q�/��v1a{J�W���]�x}NI0���ԏ�.fOe	m���h������#oM|#9���!�`�(i3N��	�Ȓme":l�nJ�a$�Y ������K�+���w�W���b�0�`
 ֢���뒒���!�`�(i3Ǒ�e}5�,���x!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j&���"�g72O!j���8
�O�@��2��.�g3Z�)V��B�1u:u����<x��u��n�G�A�FC�]s��i�~Fz��Ԥ��C�xi7�E��'Z*)�?�R��nj��P_Q����t�h��W+��W��v1a{J���&Y��V��C�xi7��U��)���Y;e�iK!���d.O.C�U��B��-V���$��b�D ML:���7|)�`�H����Qw�c4~Nr_�mS8<�n�ݚ�Н����D)���Z� ��(HJ�a$�Y dN�<@Iv��nt=:��:5A��p�$�`V1�������S�\zigzA=v)E�g�������(ӈ���m�r����١w��zj�v1a{J��湮��n��>�my$�N��o�/���;�/��@���WdM4@��_�U*�I����~uK7͍��|��W&":�ݚ�Н�K�\7}�W, D�cg�}Ņ��4&Ks�dN�<@Iv��nt=:��:5A��p[�t��#��%��g:���\��Hܞ�E�g�������(ӈ���m�r����;�x'_|~� �S���}me":l�nn��>�my$�N��o�/���;�B�'��a�/������Z� ��(H�I����~uK7͍��|��W&":�ݚ�Н�닓.�`�3BڴQ��J�a$�Y dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3���D)���Z� ��(HJ�a$�Y �C�|J3J��М�Z��N|;^�S;��k]m���r?&��AK��sC宸I))����A�m�(�QNȮ���k/��m#��}Dq�f�9��?xs}�k�����|	�WI�i�<�~�y�j�q�7�AԢ�a\蟴���P`��ʱ�O��W���]�x}NI0���ԏ�.fOe	m���h������#oM��:<��j!�`�(i3�⒍~����v�z`�!�`�(i3���o���F��+=�o$Ô���,��WdM4@��z(�ﳍ�f�_��S�>�!/�_�n�To�[
MQ9�F���"X��[�,�!���D!�`�(i3K�\7}�W,��+G��ܢN��_;���C�|J3J��М�Z�ׄ��e�S�[�k]m���E��Y�W���]�x}NI0���ԏ�.fOe	�b��r�
JB8�^C
��ݚ�Н�[�t��#��l��姹����+�Q�����zk2��|�kڲ��b�Bϱ�[��m�U/|w~S."��b�Ͻq%(���B����: ��ao.\C�k�ף�D�~n��1w{��8���/��:5A��p١w��zj�v1a{J���!<��v�Fr���IbW�P"G�wk�#�_wU|�1Ĵ��ޯi��ŁO�W���]�x}NI0���ԏ�.fOe	m���h������#oM��:<��j!�`�(i3��@�z]��C�x!�H�Z���,ߘ��o���F�������ʂ.m��K�+���w�M�7��<�1�����\�H��/Sg޶��j�}a�cf��"X��[��Q[R�7!�`�(i3�Ɔ ����;ƹ��:i����;qN��	�Ȓ�cЉ�MO`�� \)-�E��%����gr��!�`�(i3���i���w�XU'��
�:qEp�;�P�t�5fĉ>99��A0ok�׹�V���$��b�D ML:�ctj)��>#����,�ǰ?%{B��0B�tw�i�՗[�:X#x^�&����������I �P��M3�G��#'@Nw�z5�0P�ġ��x���u�Y�KG�ξ���I��RhF����u�*��?�d���&�a
�+��8n�TԁC*�o��_�Rv�䩲$��GQЌJ
��`���φ��<�6���n�4��;�jmT�#bs��2[�a��o���H�RtV�^�amf�M '%�줝v)ƍ2���l��k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��y�!�`�(i3�amf�M '	��1	�q��eԱ���:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��|I����<��}�u�?�d���&��z5�0P�'vr=c�w�N\`�a:-�I�3�BD�O�.r�r+��ސ����U��)���Y;e�iK!���d.���8-|�D���"sS<�0�zG�������&GЈH�����b�'Be���0��_�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��lb~*��s��YN
��)e�W�J��H����8�O�5���1tSjv��H�����Ɔ ���Ve��˅�>��{���M�I�h��}�~��l��-/a8!�`�(i3N��	�Ȓ�cЉ�M^�h۾�(�b�'Be�����y�?��}Dq�f������!�`�(i3N��	�Ȓ�cЉ�M�'DV���b�z'hۉ)��d�7�qĉ��%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j�_�Ƭ7~�rG[Pt�����Vx`a"�6�m��gO�J���M���HaU$kX�ڹ��/^�w?�d���&�db�\EX회�h�#5ġ��x���u�Y�KG�ξ���e�J�Pn\�pD��ZOU;��|B���r�����Ɔ �����Vd�;,���3�/�����Y_sĝ���w�R���y�U��\JD:�GI���o�+�=4V��	��yO��aQ'�����f���K�h�y�[ee[V	Q��2�P�?�r�&U���0��PW�%X�9���Ylom;�Ɔ �������4�Ք�R'cf���³5����U��+�Xa�H(�˕�Eo(d��Ylom;�Ɔ �����Vd���ة�蝌b�Bϱ��9��no �گ��h/������B�F~�o3����,�ǰ���9kn��회�h�#5�ޒ�K��6j�"Hs<�?j=Ծ���f���K�h\K�5~�k�좏1Y�����E�����A���@���~$��F��v����{�h�&T�n�2��^�5�^���������EXs70�U��)���Y;e�iK!���d.���8-|�D���"sS<�0�zG�������&G�'.�T���Bf����{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^^()��>�����U�._����P�|T����{7�H����8���O�υ���YN
��)e#j�o����B� �b��!�`�(i3���^g�6�x:�m]�c��#���F�H۷`1tSjv�!�`�(i3�T�n��aΪ�;�EIp�r~�h��ݚ�Н���w�w:�!�`�(i36�ZV	�	ҙ���˦G�K7͍��|��W&":�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�J	���/a���Q=	+�{�*&��q>�<�'���I����� ���JH����8����F)�~����H�V�n8�A�A�y���6���#¯��TG6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3�4br��n��>�my$�N��o�/���;�B�'��a�S���%�����ռt
�AԢ�a\蟟Q��ǺΕR��ӟ-�q�x�~<��w���	�e�<j��.#՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r��;�jmT�#�YN
��)e���^b�~H����8�O�5���1tSjv�!�`�(i3�YN
��)e������p�r~�h��ݚ�Н���w�w:�!�`�(i3%Q�[�J����˦G�K7͍��|��W&":�ݚ�Н�$f��_Ub�F�S�1 ��H�����4br��>�=,W�[�?�R��n}�����Hٚ�-����!�`�(i3	�)��&ghRV��R�4br���h�Һ�!�`�(i3��jVѭ@!�`�(i3	�)��&ghRV��RK7͍��|��W&":�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��#}�{��Jw��3��.�g3Zv���� )�W/πs����N�KRK���DV4�ސ���E��'Z*)�?�R��n��h
:h����t�h��W+��W��4br����'�QV[��;_��8W�w��fD�Y%ɫTK���N�KRra?��Ba�Cy}�����:�Nz�]'\gWg��	�Z�kfc�_	�Ƽ���8|bs��2[�a��o���H�RtV�^���M��2E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81tSjv��H�����8���d�W�J��H����8�(����T�x�"��XƤ5_�J�	�LÆ���#��p��;�{��!�`�(i32�#���l�
@\ه3
�v�v-}�	mp5���%�+� h�ҩ��wӨj]h���^/e��d�G�.�@��ӯ�2�`<!�`�(i3��jVѭ@!�`�(i3}�1�Ha�E�Rq���my$�N��o�/���;!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6���ޡ�m���Y�$�9����~+2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��Wv�A����w�V�"~�ӵ(r7�8� ��$d������`7�tȈ������9P�-�,�AG�<���X饿��!�iv�aQ�Ϧ�M�ኾ���L��r�U���f��/?L���u�D��D1��n������� �k,
"i�̄�ѭ���ɿ�kF��l�l"��l䋬5Kq!�`�(i3!�`�(i3}��[b:��'(K�lc���97�
C�dA��:���f���X�k�J�3���-Q�OP�}.z)y5�[՚1D$Q,�WP����jw8T�1�c�{Wo9�����<��l�Օ��qvdЧ^{�jmWᅫw�5�O�%E#P�;����<��p��b��!���?t��my$�N�����X8�#s�vS�em;����^F�=�_�7V�o��_�Rv�䩲$��GQЌJ
��`���φ��<�6��o�.�u:u����<Srƫp��xjzӝ���I(͂��-�����d�tuѼ�!���{��b+}y[�߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��la��o���H�RtV�^>�Q�c6�~nS��\z-+;X���W���b�0�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ����[7Y'��k��F$�kj�L��M����4�	��������A$�P������5d�������y�:Fa�7���W"�P�K¨}�n/�J� &�0D��xjzӝ���I(͂��-�����2��}�����3R�Ƃ�nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����V(MH��ZRR���&���Ɗ3I5=��)Q�]� ���_�hbvk~�#x��Og����1tSjv��wӨj]h��J��sr�lv{��lw	!ݞX�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�ML��M����4�	���P���/��.�g3ZE��g�Hby���=)�Vk����/x �i�{��R�S��>j���T�}ɻY~�y�����[�]9�(b���J��:����}�6�nq����P�U��)���Y;e�iK!���d.B����=1_#u���GT�A�IÙ=�H��'�PD�{y����i�q,?5q��7���9��e���W� �{Z+����"sS<�0�zG�������&G�����$ɔ9Q<ϯ)P<�ܓ�Y�B�'��a���� Ev��\��;�,�̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*_�mS8<�n�ݚ�Н�|�au�(ZԮ�g��#��ܭ i��Y�{'%sk����w�;F}���V6�!�R/\T&O���GyV�ش�oh��!�`�(i3��=m緒X�X�pF�#}�{��~v� 1��M��%�p@m�ڨ�hծ!�`�(i3��Nh�=f[��8��GM5s�FF���p&1"?�R��n}�����Hٚ�-����!�`�(i3*�9��.���=�⳿P��}Dq�f���.J7h��,?��&�)�
�k\�i��}Dq�f��߆�p�h��{$�������LQ�/8۶&��L�H�W�J��H����8�O�5���1tSjv�!�`�(i3ʬw�S���q9+t�}�ݚ�Н������y����������"��Ra])n#���r�����d�tuѼ�!���{ʬw�S������W�!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j �_�ȇLШ��+���Al+�HtB"o
�BP�@Ե5���Wd��%�o��_�Rv�䩲$��GQЌJ
��`���φ��<�6�닓.�`�3�P���F\\���F�`yx�>�+X�M?��y�!�`�(i3�4�	��3|v��Eb�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��lb~*��s�닓.�`�3p��2�H���'T���+8!��?V0D�	�I���_
�u�Y���H�hbvk~�#x�DS�AvF̓@?5�#j�o���&�2����+�+�5���4br������Ľ����Չxv��Օ��qvdЧ^{�j��@�
h����Z>ؼ��XyH�RtV�^q�\E��0�d��+��2VP��Ѣ�ʒN�ċ
�:qEp�;�P�t�5fĉ>99��A0ok�׹�m)��T<�cny��&񮣙�cq@�w�R���y����<�..�4��3�U��`�Р�(�V�'G�+R���o��_�Rv�䩲$��8��I�:Fa�7��X$_V� �6(�X)���7�癆cgQw�c4~Nr_�mS8<�ncp6Dq����Cs�q9+t�}hDJ��3��%�����q9+t�}����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н��xmQ,ۘS���VW��F��+g�ݚ�Н�ʬw�S���<v�cn@�q���uҽfĉ>99��A0ok�����F��O�\E�W��4bX$_V� �6(�X)�ҽ�6jQ����D�X��;���B�9�Q�f�����+� ��*ȑs;��|BX�D�mP�>c��?�B�t�xr�t��b���2�b=���i�WgV}Q
�Waf���� ����6�o8:4�I���c�90B3v�A���('�@�+���3f	aF�o�@OiFA� @D�H*�=bs��2[�a��o���lO	"����q�\E��0Z¥���5.�{_8�Y��=�}�Vݨ�,bxqX��k��^�1��dc�@c�����h��-�����_���`e<�Ia��la��o���lO	"�����2��}��M��V!�D�WaU��,bxqX�HN��R��bP�63Z�t�tH���]*bP�63Z�t����؊O.�x����VǪ =ա�0��L�r:|�O�E/�9��"J j�E��'Z*)�?�R��nj��P_Q����t�h��W+��W�H^��Ƨ�0͜��!?@K�,bxqX�����,�ǰ����E
��sp���m��>#e�6&	  �ιf����ZaL݊���2�"�G�p�Pڹ��/^�w?�d���&��]�o��A����\��]8��	���#�z��%]'\gWg��	�Z�kfc?�#	*]]�iI9�o«IX0F�M��ŊPTWo9���b��|2\���F�`yx�>�+X�M?��y�!�`�(i3z�
1���;%��v��!�`�(i3��������Z¥���5.�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r���s�Yls��8��GM��-����!�`�(i3z�
1���; ,��rQ�U�^)����ݚ�Н��O)�b�c�!{p85v{��lw	bo N��7�$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��o�.�u:u����<�x���ަ�I��O0Y�6j�"Hs/�n�����E�xc|�+�AR+@|#Z�1�IX0F�MV�ҁGG`5:�����+�^n=\f�5>�.F<!W���t�㮫����"sS<�0�zG�������&G��+�t2�������/��kOT�̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*�Va�ir3[�u8���m�~r�D�4�.h=�,\���P�75��iI8�ѐv2�8�n�"X��M�����)m<�3HYʨ�]�_F!�`�(i3��c��qVw���%���RAԢ�a\��?�R�_��sV�����נ2<�i������b��u��r���#�-�p����B��6�<������NM���fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx?�y�g���w�R���yxl+�����o�+��5�s�AEA�W��x�13�K��oNYzZF����9��]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7���z�G�	S�uimK������t�r$ɓǃl[�Ƶ�1tSjv� �#0xg�`�I��Wn��>�my$�N��o�/���;����������zՠ�����˦G�K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н�>��:J�E�<����i"����*ȑs��,:&�^��,Q����-����!�`�(i3R�c4!`��Bf���Q١Ӿ�$���l�K�F���m¡HN��R��bP�63Z�ta�F�������Y���D��3��bt�u�&��F�ߏ��D厺��+�̟�1�8�>r&�G�p�PPS�H�I��I0���ԏ�.fOe	�S�4��=ǚ�-����!�`�(i3Y�)�}��EXs70:���&�����|�b���Fa>t
�:qEp'{w#/ B�d�tu����a{���Bf����{_8�Y��=�}�Vݨ��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍʞ3���h��[��1聦Ά1��<����i"��@#('�cH1��<9Oy��]#�0D�	�I���_
�u�_C�7�2������}0n�V2���]#��t�ѕ1��ŦL�ݚ�Н�!�`�(i3!�`�(i3'����t�Gf��x��9	4��t�f��x���<d3"������-ќv0D�	�I���_
�u�����|�G�p�P��<jV���\�H��/Sg�w��'o�+u�d��D厺��+w���	�e���0��Qܓ'{w#/ B!�`�(i3��7I���|ag��6��+jq����i��gE��[4ҹXH�m�w���i���Z���D�U�2Y��i�p��+˞j��&����Q]� _ό���.�@?d�s�8KFmғO�4}~n���,a�n`5�fK�\w��0]\o�LCd��.ZQ�*�3���g�7s�9���o>��l%i�-}�
�?���B@��������/s9�d�٣��>����C�b!��u�<�`A��_i3i 
�c��]�!����M[��ǢHe�-�c��3E M0�F�T��BZ鎬�����	�7 �#�E �����	(��7�зq8�Ј'���Xw�j�7����w�K�b��2W hbvk~�#x ��M��.ᬵy��"C�����T�\ �͹g}|�H�I��'�!͙��04nԴ�V����U� ���_tE��gVB�3?�J	QT��8&���I�%A?�dL+jq����M~�̀R��n	l��Q;�im��ȍry��	.�n^y���\+��R�4.����P}�=l�q�������g2��Ɏ�#���?�5q{! l��2
L./;�Ly�Af�?ǉ�=�e�MW��Rj�q�wxo�~]�g���[��}��#J*�Rs�08�b(������l__���#���,Wc��I��@�hGq6��nX��U�	vn����R�����_���!�`�(i3#B��F�!�`�(i3!�`�(i3��*�{6��(�w���!�`�(i3Y�"O���j����I~!�`�(i3	�=��G���v�8:ۛ@W:���#���F��n3p_�#2\z��o t�J�PM�Y��G%�&8�,�H*W��u�a�ݚ�Н��^yE⛀B��+ H!�`�(i3ˮF���t�F+������X:��+�i�	��_�V!�`�(i3-��w¹��<d�,��L��#2\z��}�� �с�'(�U�c�&8�,��
�Q!}-[BvGޣkQ�A���ۖ$����nQ�rV,?�����ݚ�Н��V��(��sW��|E�q��w\F��G8T�w�nf�?ǉ�=���S���_�������"�9(���l ��ǣ©���u��4��#�N�X�!�`�(i3�M����iٛ[�Z�Z������s��+qѭ�+g[�</Sn��-�¾L��8�$��`���VF�˷�f�?ǉ�=	s(D��&8�,������	�;�ݚ�Н�4?s����k-����b=�`
 ֢��-�¾L��8�$��`�� ��M�#f�?ǉ�=�ϋ�LΗO�&8�,��@��Y��;�ݚ�Н�*��^�"~H�҂��hWj���H�D���dݮ%*!�`�(i3���_͏��X;p`�����G9L�bW�mT(�l\�6�'����7Z��czZ����N��E�Es!�`�(i3��w]��&��)��>.$5<�`A��_iN��E�Es!�`�(i3)�{� �"�X;p`���2�b=��<�ry^���i�\!�`�(i3�$�~c/v��&EA)<�!�d�<�-�����q$��7�H+�����s��߀������k-�-�����@:[�X�	�J�`Ԡ��`��!�`�(i3��	&�K��2q��'X�qp�c� &��GE<�!�`�(i3�U�s
ƺ�+e;��5&�(�R|�G᭞���Np9�A(jgOR��/�q#a�_�̞��>��3
�v�v-}�	mp,��_А#�<om�����M��2;0��L�r:�9]��j�W>l��? Ah�*h,ChW+x⣗�C��ҷ�㗼�?�S���J8����E^��o۪��5/:�� N
�������?;����IX0F�MV�ҁGG`5:�����+�^n=\f�5>�.F<!W���t�㮫����"sS<�0�zG�������&G��+�t2�������/��kOT�̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l����� �'����u��r���#�-�p����B��6�<�������G9L�M�7��<�M�l��S�J*�Rs�08�b(������l__��E� )�&9*�����fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx.F<!W��Y���x�wbk�$ *�������U��RbAvx��բS��\P0RP���50f
V��.ᬵy����� ��g H�8��#eW���Z��1���~!�`�(i3V[B�5�mw�R���y>��yС}������Rr����t70�6�H