��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω� C�`N��D���ÿ0�^��p*z�w4G� ������[���a�8%`��4�s�6�XAoeu��a@����þ�V���	��U0�4B��A_�1�:�Ω� C�`N��D���ÿ0�^��p*z�w4G�� ��d�n}K-J��K��z������3�z�ω���D���+�	���lF72��{L�8br�.�/�d�������4�;(�GoAW�~.8%D.��n�P��<2�q�U��k�8u[\E���@N1�w�0XL����[fe�Hs��9lSUQ�S��)���2Ee�Y�R2
�I.��	���
����k�������0�?�}4��ѕ�������U��=>bMab�	;4��G����a�����(�I�?g�f��r�F�5��I^ξ��ݴg��S�ZC�L|�w.j��6��H4�
� �AH���g���	r��ܤ���=���Z炈\a�T�F@�4%�����^)�D���%�d��C��m����߼��:h�I�?g�f����~����/x��-w}Úl�� �'m����_m��+++�i'��Cx�"T4�^�o�M��Yј���m�!=�y����h�}�_nR�� ��/��OY�N���o?�M��;]�Xa�v�Q�W�%-C��oW9{:n���;u���7�r��b}()pxt4���J4xʆ�7���I�9���1� c��(�U����	x]�<���e�P����>�]!�ՄN�Ӿ��)�$�����PГ��0�w&��EO�{�������E��sޜ��*�c�N!ͬ鏈wƠ��ѹ?�����qU�%��Sr�'hJ�.;��L�OT�+?3�l� c��(�U����	x]�����O���8�t	;N���=��B�3ʦU�:�%�+M��m}on���b='��\�4�sW c`k��TT	q��$f��Z��FUR�.�;�~�MUs �ˠ{�t!�.�r�c^�e���zǒBs�&���b�!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�
+&�s�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v�lf)@̲#;���(�s�-���f�i\􁗊�n��\v;V[���b�/r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[n�+�Uz�QL�W*g;X~09h�i��I�?g�f�$��P���o[��+��T��٤�2[51g~Ӝ��ajƎ�c��(r���U�2�C�b��}Y���%�5�1�:�Ω��
�/�r}|��ι%9��oGo�Z�J��ݪ���AOge�����Ӿ���	���q��q�©������5X�/x��-w}�USֈ�����M:��;6aJVlO/8֩]=$���GZ>.�0�[7�d|���XP����
/1�&��F�r�f�teE(��o���&��J�1�KB|1<\�ԌY&�xL����J?��\�vňu�,�s���2��̪U��֜��3�a�\����9�	��%�t�&_���9� ���3�ҺIÙ=�H�x���������CgU��d#]=�~�n8M���dbP3z}�&��ٙ���O����
�}�=Ll�����,۽���}i�@�5�}�]���=]A��O�T=�4e=��-�ĕ|G���c��� �G�T(���D	��U�l>o��|�l�n3؍��R��j�.(Wx*���Mڷ�21!t*x�S��|g�Y�'���Xw s4S�'�i��`�z��GZ>.�0a�3�9�nj�0��E|�,�CyW�f�tR�wX��q�\E��0	ozqP�����
L'���Xw s4S�'�i��`�z��GZ>.�0T$��V�������CyW�f�tR�wX�����?�N�By3��<Z鎬�����X���*_��(֥�S�)37J*u>����CΫa������<��z��}���w�V�"ev�mS��0�-����#u��Yk"1/|sL'���oֲ󄰊�
~�d�9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6ea�8���B����g��Tݭ�EB�.���mtL�iײ`��I��'��۟b�/O�=�ͦ����Jg�Z�n��[���M��Ҁ��@F�O��eτ�bs��z�h��4h���}둮c_����+�˂߮<uMՙqL�m��0��E|�,�h�p�x�������c�A�L'��!�a��5�%]���a(􆿳��?ƾ��,�&� �L��ۊ��|����OxtX+�Y��M��ҹf�f3'����V8Joh���}둮/��q�&���N����]�u�L��ۊ����]��i�"�`�|��K�z��|����=%+]Bo�A;h�F��O�i���AԢ�a\�P����ˮ��lC��U�T�\ ��y�.�`L�P7koеI͢'�����t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s��.|Z���I7��-5��6��	���`y����@����gG��l��`��y����~G��a\Y���{lGD�V�B��иܖ��A�.u�r���,D�=P��[#֫��/f��Ԝ�]����n�4�{lGD�V�B��иܖ��A�.u�rI����"�*�şxˏ1"Ohƪڈm�d�٣��c�A�L'R�o�����5�%]���a(􆿳���2����.��DP֞ �(nyfW��􇃬Tk�H@H�֦g�㎏qló��@d���/��=��K�R�hE!3��
iEE�G��V �-���W|�M��3�j��gGD@�F��qt�N$	L݃g{~�5��'x��}v�Kv�LM +�gf�����w]cH>��DN2��J��_1��'n�^0o��S��S�B
��aP/;D���Y�������eŞ%�ޚe���|^�a�u@�3�Y	��
�t	���+�+3�ϡ��]Y�� ���9��cKԾ	I����`�z��GZ>.�0�i�ܰAe�0
A���̹U�����r���	w	Qrk)�7JS�����,MLG򬉢��S��ȍry��	��yso6L�4��'��v��@�������>[HÛON�?��!�`�(i3,ԯ���gn��Ab�%^��}Dq�f��N�v�1�c����L�{�E����F�Z�>)�ώ�~+�ݗ�r'Z1p8��e�j�!�`�(i3,ԯ���gn�J����� ��}Dq�f��.��Ԕ�	���ZX�E����F���8�TP��IL;��$��8_�8���&�'�al��p�I�PD�na"�,�>E��4];ˍH����TI��Ԫ,щ�"��Wʁ�Wp7�:�!�`�(i3x�]�V���t�����[F�a�+�ީ�%��Wp7�:�!�`�(i37�ܥ��2�`e7��9��×�>���`�)J*~���f��0�5tU���D	��U�l>o��|���bǬ�=��I(�c��U��j�fH��>d]=]A��O�T=�4e=��-Y�VN�=��7p�J��PWV����ft���}�k�����5	��{�OF8F���m¡�����hWK{m35%7� ��yDgx�]�V���t���CՐ3��F<Y��j3��� Q�N��*���������@�%�I=�4e=��-V�׍A�ž_�F���yso6L%+�&��v��@�������>[HNl����!�`�(i3�E����F�Z�>)�ώ�~+�ݗ����>[H����&?�!�`�(i3�E����F�Z�>)�ώ�~+�ݗ�r'Z1p8��Y"H���!�`�(i3�E����F�Z�>)�����˟y� �>��|���;��x��B5��E����F���8�TPm=_g}b��t��6�5�p���PF��W�!�`�(i3зq8�Ј)w�<�_N��M��+?���C&����Wʁ�w�*�fBg�!�`�(i3���+�J��U<o^.K�}�{��$&XT
��"{phDJ��3Y� 2��4����7
!�`�(i37�ܥ��2�`e7��9��×�>��� �>��|~���f�A�������E����F���8�TP��@E�`�8���&�Q�$_��^�|n�M�!�`�(i3=]A��O�T=�4e=��-"w߻Y��}Dq�f���R�㺺|:=�C��Z��N�l������l>o��|���JLm|�Q'݀�=���SCh��{<qH�~�!�`�(i37�ܥ��2���kܪ���*�LNm�t����}ꇐ�622���k˗S�d�!�`�(i3x�]�V���t�����[F�a�+����ܗ�J���z!����k˗S�d�зq8�Ј)w�<�_N`E�cvR+��}Dq�f��v1a{J��]��3a��!�`�(i3���D	��U�l>o��|���bǬ�=��I(�c��U��j��k˗S�d�"�,�>E��4];ˍH����TI��Ԫ,щ�"��<H��(����O��B�r�������5	��{�OF8F���m¡�����hWK{m35%,�!�H<Ȳ��+�J��U<o^.K�}qW8+����8���&�qr�^*4y-X��;^��J1!be�=]A��O�T=�4e=��-V�׍A���}Dq�f���*����	��Y��71{!�`�(i3���D	��U�l>o��|��b��7u�� л�b����\�TfZ!4Я\�rƛ�}�ٸW�{vK &�k+���!�`�(i3!�`�(i3=]A��O�T=�4e=��-�z�)lq���a���8���&�1籢��N�o!�`�(i3!�`�(i3�����5	��{�OF8�_�/�ߥ$Nx���t��y(�����������(������%�G"QL�)w�<�_N�eب�-�t���k��-��Wf<��;����7�/>�"�Ax!�`�(i3!�`�(i3x�]�V��;���Ӧ��Gjh�rO-�����`J�^���gJ!�`�(i3!�`�(i3�E����F���8�TPT֟��B�:УWKŃ����`J�*���u�Ww3i�|�!�`�(i3�E����F���8�TPT֟��B�:УWKŃz�q�����GO����!�`�(i3!�`�(i3�E����F�Z�>)�����˟y�u3v��U�DnK�]_!C6%K�pıN�c뵣�"�,�>E��4];ˍH�,t����t�&Fc$�n}��]"danS����˥����AB9���w�!�`�(i3x�]�V���T�3�R��	���I����r����$^�y1�\GD@�F��qW��Ґ�Yj���|��1��$�V��b�s������=���aI���;E�@%���8�a�"��FX1��t��L̿��$|�/|�z)�_m-�oq��f�}������!H�P|�����7JS�����,MLG�	�6���I!�oLS�)37J*u���{��}!�`�(i3!�`�(i3!�`�(i3���w�P���+��o�.o�`��K5�w,��"�����q��l0\4L$ֵ����門�ҋX����Q��C� ��!�`�(i3!�`�(i3!�`�(i3k��j �%��:wJ~��r�=��uy������I �P2<WV��
i�c�rד��L��T7Ê7�E�4'���Xw!�`�(i3!�`�(i3!�`�(i3!�`�(i3 ��ii����1��뜙��L`Q�
_�J�g�J�LQ��wEOJ�uxm�!�oLS�)37J*uc�A�L'�t�Otj{%��ߛ�8���/��}�Ш���my$�N��;� ��b�� л�<Ct�a��\=��
i�c�r�]���,q�7Ê7�E�4'���Xw�j�7��k�-i�9~�,0=]^	�&�e A7YzE�ˇ�h����2�[Q	��
�Q�}#�ҒIs{JE���=���B�NoSƏw0���|��*��<��z��}�0z�cUL��լ[po���̛i���7�v�ԯ��Q[R�7�Mei|�{LZn�+�m�&(|dPSM0.�J�a3mPy���dn����]�!��	Ǹ�y85�&�;���
��#E�>���T�\ �͘�f��p�b�z'hۉ)[텡#����Mei|�B��Vj��m�&(|dP`�,����}];�SS<-S�N;��0�"� ��w� 9_�똣w�ٽv�yq�`0�|(O��"��"�T�>�#�ҒIs{�D������:_�_5:��(�I>�IP�b������:�kR�$fOyQ��������b^��ɮ�� л�G/1avQ�e�b�����,��Z?m��r�գ��(W�{fy}P��B�wo��<�,R�8Ġ��x�6Y�nlH�I<�6�Q=���x��<�6�Q=	I%Mq��`Ҧ�׶!z1��,,ҹ�$�OD��G͘B./�<ĩ�46�;:��/k3gS�yy�ã��&�զ2p�$�W��	]�	���F���X:����*�`��g>~qA��@����M�P�;���=����t��LӰ�+M�ҋX����L$�����/���NM����s�٩�삂��!O@T'���Xw�����U�VA�ڦ�c4G��.���"������O�69:�BF�!���q�%��Ro�����:,:��G��.��M�zp�p+!�`�(i3!�`�(i3�ܒ.���T_�[�S{�o%^�G@�m�񈽢d@ǚ��ظ���K����^W��k����I�!�`�(i3!�`�(i3�Ѳ��aS�!-�+_����1�"`��Ę*��7��S�S�yy����9K��r|Z�%%�5�_Z鎬����=���ޒC>��}Dq�f�B)vظ�u��o��C!T*p�VU��Jp��T���ȓM�Me��d	�A��7j�!󊾵�e�;Pq]g\ ���ǋҠ7�	�ߥ�H�^ /m�6���<�6�Q=���Ң�Q<�6�Q=	I%Mq��`Ҧ�׶!z1��,�У��a�p���L1�%�1��zo%M|�e אN�ʡV�l��� л�G/1avQ�e�b�����,��Z?m��`�������VRj8�@��"�VGN�Ar��$x�y�ˏgԊ���c�.D�#�ҒIs{�>Y��}�:_�_5:��(�I>�IP�b�����LQo������R��H�O��	�d[��K�pHj�4�\��F���77AƐ^�8�tn�+�e��j�3����&Y��V�贅���Ǯ0��]㯟B./�<ĩku��j�,�J�2��s] U���v{:��h��MB��V<��z��}�<ͧ�:|��b+}y[�MQNv�2���!O@T'���Xw�����C�VA�ڦ�c4�5Nleo���_�n�<��z��}�<ͧ�:|��b+}y[|�\m���SLq�N���])���/�Z鎬����Ĺ#{��ž_�Fȼ�Ŷ;���@��O���Z鎬�������(��變�\_(����O�e��3T{�8���/�l|�*"k���(ӈ��4��S;UA7��I+��ė�?�����m���B�No��I(�c�]C�:���<��z��}�0z�cUL�k�	����V����fta�ʱ�RK�7�v�ԯ����fbK7͍��ճ��)�ȓM�Me���섫�So#����a�kEӮY�E�7L�V�wļ�T���
(dP|�����7JS�����,MLG���;EF����TD���rs�i���YN���G����exa(􆿳��_�"ۆ�$�D5�bY[r��  G�E
b�+|�����
L'���Xw�j�7��k�-i�9~�,0=]^	�&�e A7YzEF�d����:p�NgO<���O��ڻC�i�e�0
A�����T�-���.�U2@f�Û��ƫg�T6����Q�u;��|B�]Z#���ҫ��N�-�R'cf���³5��&l�����#W�U��ظ�d���!i��������7�,��n6�o8:4�I���c�90B3v�A��d�G}%����3f-��cR�O�wFlE� ��\���F�`yx�>�+X�M?��y�!�`�(i3���_��������صW�my$�N��o�/���;
�:qEpk+Q�h'�Ȝx�5W ��̫(� h�ҩ��H�����Yu�������&G!�`�(i3{k�h�+�QCj�4ZP-�O���7�:5A��pfĉ>99��A0ok��fĉ>99��A0ok��W?�;���^�#�n=��ht��HN��R��?�d���&��"��aT��3G?�d���&�Q١Ӿ�$Mu��G�ا��а=��F�5(��j���rz��Se�������,(%�����Ε3��"��;_��8W�w��fDSbp}���y)蜶��3v�q�ٙ���O�Dw
�
�{��_r�e~��:�5}`�&ڣ �#A=�Љ������qθ���6j|ݎ��;_��8W�w��fDK��lG�?"���\�)��E�d�-���geW���w>��Y��d���!i�^Xe���:��j�3;R�Zם�³5��&l�����#W�U�����$1&O�����%kR������ ��0���u%?gV��U�x�l��1:�N�*�x\�
�=ĭ,Ϸ�@��;!�`�(i3��4��#o�;���[�����&��[&��YF�"�����G�ݭ�,��#Ay������|�vh_n�,��v#��At�B7Ԅ����$_��f3��"�2VPڢ7���w�E�V{�!�`�(i3߼��� �x� ]
� �SI�����+6�l�?�Ho2����q��3[�[�6Z��et<� ).�xz�\�{<�?�Ho2��2�n������Ir:�fC��T����ܼޥ0D���>M�J<0L�J��2����`x�dˆ�ָ�K L��ݚ�Н�K�± ���.]̌�+k��eژ���Q��K�&�C�/¥�����Ј��wf-��w¹��<d�,��L��!�`�(i3I:�K�R����4�txj����R��á�~O��7�I0I/R�R�)d
ӳ,\ͨ܉p����O,8�ݚ�Н�P�I��"ĳN>�`������	�;�ݚ�Н��6�5�p��`�T1)��/Z鎬�������(���G�n봈2=��At����G�̝�hy�t�]�|����*[UxG!�`�(i3��9K��r|4�:���m�
��,!�2��}��g��9|P�wAA�Ɓ=��2�[Q`��l�\m�(�:�f,�c����L�{��n�T���#�-eɤ,-L�	�.���ǖ�!}�	76�&�;��|Bi��_�槴��;_��8W�w��fD�8qlL`i��v�%�zq_҂T�q�w��/��=��K�E��{#6�a?�d���&��D�U�2Y�e��y���vWދ�qc:P����ˮ�����v�h�g��U-�e a⣃_B7�}�!��K�\7}�W,`q���9�z �VBD�!獜t�����Oxk*����.�g3ZrZ�0m�\�S��u���.�g3ZE��g�Hb麭�H�κ'��G3#uV��rU�w�⽒��8�>r&�,�Aٺ�H�f>x�:	�W+��W��?��+�|EYzȧԡ�/$a��F˯�+)�+#c����nS�3�ǻ��d���!i?V��j�c�N�4��@Dx?IJ��a��L�x��5��.�g3ZrZ�0m�\�w�|J����;_��8W�w��fD�W�_�����!b�*���VU�簦D�L�x8�̹�y3����&=)X���37�˱�5�6i��̨D�:ʽ�f��q�	%�t�B�6cڥ9��[���"��Y�Q�qF`?3S��n��@IE�U����S8��y�)xʔ���V�� �\�HP@�a�?�������o��C!T*�q���U���0��t��!��� ��]�!���/lwb���&�v�x�o��C!T*Y�{'%s�Ǹ2���_�A.��XU�Q�*�g��U-�e㩙�#nr��⹌y��o��C!T*Y�{'%s�Ǹ2���_�A.��vV�v��g��U-�ewǓ��}�K�bO\�Rэ�ҋX����;�ƀ�'͚+�0\�N��{l�f|��rs�i��s�٭��?��?��T�\ ���-#kt�۫gwD������m�ep��Ve+&�&37�˱�56,x.���G�9Ҥ+��o��s4k�r�j�b#���xf36�x8@�*�p�ɹ��I�``%|5��0@���&���� ��
fC��T��9���!�a�+�wVi�W�W��<��W{0`ꄳq�Y�
p�-�L�~���A�U� ���_Y�VN�=���M^���B!.��@h�^fC��T���	�5IW���-��v�r��Rϻt<� ).�xg�"z�JmD�?�Y0�
��аJ@o�C���j�}�X��>�SS�]si�O�����rRV��F��s-"&6��\���,}	f��ņ�}h$�q�BZS[]��7^�� T��,}	f��ņ�}h$�|�7����s�ݺᣄ2m>y�H����,}	f��J�/`0�����������}�(C#ƀ��=���a��JLm|��� ��,���ƸL��؅��FJ��o�C���j}�<��{�gؓ��')4];ˍH�� �d�Z[���0�2q���=YU�pSVL��˚�'n�^0o��H�3+ql��緺4v�r��Rϻx�]�V��v��K.Ū��lEs�l��緺4?s�_{X4x�]�V�����TI����G<�̂{����Ka�Ġ"\R؅��FJ���d	c�b���� B��lfR	�_�]_�9M��v�ɢ������=���a�`��	4Ij]�������K70y�=`HV7�ܥ��2�/��:M/�V���k�=��`
^8L���o��x�R5�A�yx�]�V���E�(��� �M������勤U�N�"1��`&X/64];ˍH�O������=򩦞iQ]pV�����ٙ�����\�}��n�4];ˍH�T֟��BП�� �ׇӭ��o64d�kʔ��>һA.e�@H��F��5������'!�`�(i3!�`�(i37�ܥ��2�`���{�L���i������Fz�z��?�F�ʙ��9���!�`�(i3!�`�(i3�Q�^�y�zL͊�q�����7�f�ޥ0D���>M�J<0L�J��2���!�`�(i3!�`�(i3l0��F��j �i7�sp>�(��&��^*?�z�̒�7�dz�H!�`�(i3!�`�(i3"�,�>E����\�v�Q�x���sȸ�"rR��n�1����]���!�`�(i3!�`�(i3���+�J��U<o^.K�}�d	c�b�p��I�=����d�|���=�Ҹ�S��F��u2�k������U<W�L�x�]�V���n:�t�c{DJX</���m}����뺨���¥������c�4��s���rۺ�!�`�(i3!�`�(i3JHn��z���G7�����Fz�����$G���?E/6}�U��!�`�(i3�Q�^�y�zL͊�q��r{= { _}��*�