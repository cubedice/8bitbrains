��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��U��}��x�� �� ������[���a�8%`��4�s�6�XAoeu��a@����þ�V��1�Wqlw��9�K���m��+o���sp%��X�����b1Ø^���#K���lӧIA�a�V��R�z �:�؛��px�~�J�'�دv)h�V~�$v�p��"}�v\-8�����Ȫl�M6�a��rl�ʩ{�Bfळ��)���X�$� ���jǎX������n�q��}�p� �Ñ�]�*�p�㈍x�!����Y�f��a�Z��Vb$���N[E�=����tL��	Z�G�a}CK�fC���4�O�"�F�È���_�O��<$e|����w'��1�:�Ω��U��}��x�� �� ���������	x]̢/����wЯ�mڍ'T����X�w{������:�%�+T%2q򋙔�M-US-�8<�n�У�Ǝ!�ѠV�>!�/�7��u���nEA��x�!ԝ�{��/Ƽ���\�4�smg�:�TZz�y$h��ݔf5*`]�|$ɋ��c�~�MUs c�+պNE��#Y��#p��'��������S�����:�֣I���Y/��S"�:����:�wl B����/��;��|B�6L����k�y.�)$����\�4�sc�[�.����xy�V�
7w��C��LzX�AX�~�MUs �.Eٓ�9PHvE�	��5j�rO�r�O��C��0��ùh���T�mߍu�M9F�*AJU��qχ�V���7C��H�j�?`%T=1�)�f�0��H��k3��Ԩr5@��_k���f0� �B͛	�m�O�����<�LZf4Q�����RL�a)�ƞ��U<�K�?g�W!ǫZ�<�F�Lo��i'�7C��HM|C`r�3<0��:�.u��w)�S�5� �7��Mv�9*���f��^(��f�)y�8�:r&@��=��$얃�rb2 �Q[1I�����w'�\�Q�3M���e�t��yn�	� �x�m��n~�q({L�51��;����'��%Ճ�86���H�aF��6��I���j�r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�E�s��bc�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i��I�?g�f{*n/�,傴����'SR����.�}|��ι%9M��j@�����nEAJ_�'��P9��3g�ݜ��s8[Z�`
5��*�zM�D_���.���nEAJ_�'��P9�tw:g+��T��٤�2[51g.� -��E�I�?g�f�$��P�`
5��*�z��Yk"1/���%	v3����M�sKJ�lق�����'Sea�8����g��J'�{g�P�r�|Aڙ���M�磋��w.V&��B֥�(����5�Z��f��Ո��D��2E�uq9����ea�;y� ����t��w¹��<d���<
DN�%Ah�%4
>��XP����q����}h�5,Wlr�r%)cA��u*K6HT�����N�[MD|��Ld��g�U��֜��3JHn��z�_c)���8ӋL�o'hnuZ�v|��.���hGD@�F��q��W��I<��fҾ��9��ЂDa��(O�J,����]�!����M[��Ǣۧ2���{��j��\w��0]�\�LtF���|g�Y�'���Xw}T���y~:���_L䦅�{ZC�$j'���Xw�4��}�<ܣ�<L�|��]���c�A�L'��!�a��5�%]���a(􆿳����^���`��׊���TD���rs�i��d�	�6%Ld��g��5�%]���a(􆿳�ؖ��d�I�� �:&��I�?g�f�,�� zr����$l-�㰻��������Ls�F�%ܪ���PL~΄gO�3f��*����"�Q:�{�1��q�©����y,�m��M�5���9���$1m}�
�?�����}���=�?I��)^�q�bx?������lC��U�T�\ ��i3�|)sՀ�T:���V�s��ҟ�s�_E��V�no#��٠R�^Ƒ����"X��[��Q[R�7����n9�yE,~��7s�9���o��S8��Ѽm����x?������lC��U�T�\ ���>�����+�@��ZZ¥���5.>�W��*(��F���5�L�1p/-��P �R�)R7x?���Ա��E���2W���R0�����wc�!{p85c1s�B�~�yӮ�)��	n�1tnzʘۥ<3�\"H��E��F*�L��!�`�(i3�2��}��+�n�)����%�!'G�+R���o��_�Rv�䩲$����x|e�Fd�G}%�ȏ�%|������"sS<�0�zG��� ߛ��u�����j�Bp��vdN�<@Iv��nt=:�v��؄aX���$���͜P_�_S:g�RMm�o��'����d����3�H�����Yu��� ߛ��usȸ�"rR�+?B�OA&k@C�Ɨ0z�cULb���H��u:/�ˇׇӭ�����F��O���uZL��\z>�L���$H��)��os�鮊W;§`����;8Qܓ<bm��+�Z����y�+��Y����S���� "5�]¥������]n��-��AE�HÇG�ݪ�򈟗��6%�a�����ݱ��������l���Y~�y����6d�dG�7:����b���4��)+�[Z��?d��A �4<��!I�aJ �!,$��:�e�hfH'��!�i����VZDf�?ǉ�=�2*Q=F���q/���<�����7
��+qѭ�+g[��_F�k-��苇��Fe#OOJd֯̇i�d�?�4�0 L?�p���@Z��9��稕�a�/!O�f�?ǉ�=扈�0��"��S8��@2A^=w��;f-�2��}���zgm##��+?B�OAZ��| �Ɛe�v��ҵl�]�!��	Ǹ�y85�r5��=m+y�-\֐��k��m6[��-�b�+�