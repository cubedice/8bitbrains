��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}����M7\F���r����&$9g8�M>PFWD#�z":���ӳ��_�x�$t�`a\�R�F*}Ø���K�ZF��W��`k�ZV"���:��#tC������s��n�
8JA*z�w4G�� ��d�n}K-J��K��z������3�z�ω���D���+�	���lF72��{L�8br�.�/�d�������4�;(�GoAW�~.8%D.��n�P��<���-ZW�tZ�+��[h����jǎX������n�q���xP����_�L�P�:Zqyf�F��'�Ə���ÈD6�\꾄���x�L�:>�	�$[ExI+r�� 0�D�A�f�mX�����j.�n���d�kⲽ0ۉ�@�#m��̰]`����}F��֨f,��S��f0� ����D��IG�"����[�eF�70��D8�(b�����J�E{F!��,���v�Z*���k� �\1^O�;�|���"!���5�Nn,���J��r/Zw����tq��jC\�R�F*}!����P�>s"�Xu�=�kM4v/���b��Nmj�V��v�m��Z��(Fn{�^l��R >��?	aR�}�����|�Enz��o/S)�ns)��E�$�H�T�.�P�-c��)\��A'�M8�JȦ/1�ɦ��fD��K��:�Uu�5��i	kT
�E�����l�����M�TRucDY��9�HϿ3c5M:�`�v�Uʮ�V(Y������e�(Ty@�Y#��yl7�	�=5�5s%6�%Ë"*�����Z�+�vF�ܓH�;G 6��M����iN_�c4h�C
)�R2������P��3�b����f:�_�2nW��r��� v�~D�S8a�bY�3�E��'3�*�������&�?��	м����\�W!I۾��!&O��r�����L�Y�=�B���sR۹"z�-�#�eQs�$ʧ�x��6���jm'�-��9�'���4��0:���Z��_"�q��;�8��sd�`W W��0H	�m���E��ޙv�	�"x�����
	jO��l�<u�#�$IX�2��Qb aЙ�/
߮�����q	���ޥ�i�F46���S��
j����;�]?��'(��>!XM�#�����0��G${��0�4��Z���ʶ�Z�I�"�7�\3��u�#�$IX�_r��--Sa�Qj���;�]?7#1=��*�WvO�$n������42,ߏt�}�oQ� ��紕�>&S�XQ���pU2j�k��+jGpJs��}]I+k�-�0��,��u�#�$IX΄,�H'u$ c��(�U��_�4���T%~ɸky
{:�#��Hl�P��'��Ad�Sz��=k� �@�����������ze�@!d��=���(R\֎u��·i��RZ�q�PO4ꛤ).�޽��g�7Ѝo�}a�C�|�[]?=�=\�cZ�Џ��"k@:G�4\�8�/n�G���[%y`O��@�f=H�����;�B�|�[뙴�=�u(j:�mſ���S���*�`v�J�#������g�q��5&��=����7Î�uP�T�U��%a<��A�7��m����Q�yIy{~��L>6ϲ�Ϝ���}��FB�0�sX�9���;q�j�B�C�*����%$�t� Z��i���ȆE�GVn��Bw �ͪ�(:�J�{|Tl�@�7C%��ـ��f�L�1�k�mA�����FNIR���i+vZ{w�c[��m��q6�B�9�')�J_�
W/7�䬢m]�fB�f1I�����w'�\�Q�3M���e�t��yn�	� �x�m��n~�q({L�51��;����'��%Ճ�86���H�aF��6��I���j�r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�E�s��bc�Ѽ?��Q2�=W�֯�^��N�&��^˻f��sKJ�l�i��p�7��Z鎬����@�Q�2��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i��I�?g�f{*n/�,傴����'SR����.�}|��ι%9M��j@�����nEAJ_�'��P9��'p�@�I�?g�f���\X�<����8��UWJ��)-C:����1}Kط��4�=�� F:��+���������i��i3<�f�D���X���`��wl��h��"u����i��؞�JHn��z���z�O҈�u�;Mjq2r0b�waD�����Ặ��Ϊ�Q� ~���]�a�=L[|��o\U|~'��q�S<IÙ=�H*.�PS�����z7�Qu�	�'T8�	A( ����_�h3��{I�Y`��\H�WI~�Ct���?�!�`�(i3"�,�>E����-��%Mό���.���|��p�G	kp^y�E����F��j��\w��0]�+���42�����Vc6�
f�L�qzʕ�a�N\�����ꢤ�Ogc����L�{"�,�>E����-��%M�rs�i�نW0��;�¬pX��g��U-�e�,���6+��c�r%�1�#��d_v�ј�"��Z鎬�������(���L k#Z�.T�J�� m���"u������A��o	�g��U-�ee�@Rv����my$�N��o�/���;(@X~�H:��1�, ��C�]X�.we.��xu	�>��l%i�-_ve����^́|�A�����5	���]���>����C��(R\֎u�⍽аYl���#�]�!����M[��Ǣ�J�g�*��/�p,v�ј�"��Z鎬�������(���]�����|#9���+���42�����Vcع�'����3z��ϟ�]د[9k!����N�1�Ð
�%�э�.g"}�p����|g�Y�'���Xw�.aX�bAKj�V��v+���G����(�
t�ژq���U���V9{)�7�]X]���������TD���rs�i�نW0��;�¬pX��g��U-�e�,���6+��\�2��s�ώ ���]q|���(Z鎬�������(���L k#Z�.T�J�� m���"u������A��o	�g��U-�e�,���6+��\�2��s�RdE�̈́|�]2�y�Z鎬�������(���]�����|#9���T#�3�["���'(�򑁹��E��@IE�U��>��l%i�-��+g^l�:�NI+���"B��$I��w��,�񁫴}2��8X���4bS�N1�	(f�`��2&+��T���jB�Fg�Y씤`��p]�=�_ZQ㢷F}�#Wa�b����y�E�nwE��S��}|��XH�����,>$+W��� j/~.)��3\�R�F*}�c}��uO��������uq9���
iEE�G�U�W
8�{<�����=�א=ͼ�\�v��\aьIR=���|�F(��x���hh�����RY��1|�!��3��(�����Åo{��l���h����V�@M�~���������X�7zs�p�rga�8h�Z(.V���w�c��l�,�B��+ Hxg`�H�4��`t�A~�@����gG=%� g�Vv��{
BjU-j�`�U���q�
��������n9의�z��l dG�B3�����Q]� _ό���.�}�
�?�;�j���Ѐ�K��зq8�Ј'���Xw���,DU�m#j[�M����"�,�>E���]�!����w�Հ��Fr���A�qIp��K�ڶ|e��7s�9���o>��l%i�-��B�D�F �%�э�X6و�cµ�Jn,���`�rs�i���Ӧ�am�T�\ ������q�f@�>Vۉ�!�K�&�a�M����*�7s�9���o>��l%i�-��B�D�F �%�э����y����Q]� _ό���.�}�
�?�x�j؀O��(�\G�@�L)r����'���Xw���,D�v)5�Fo�7#1=��*_kV\�헌�]�!����w�Հ�>Vۉ�!����0��G�|G�N.�N7s�9���o>��l%i�-��B�D�F �%�э��5)��Z^��Q]� _ό���.�}�
�?��(R\֎u�=7�7K�PZ.��0�W'���Xw���,D�H�p0�����dܟz-�;�g��]�!����w�Հ�(.V��������lް�l��7s�9���o>��l%i�-d�x� �qC��|���8�{�������Q]� _ό���.Ӹ@����gG1N����F�1�#��d_!�`�(i3�n`5�fK��0z�cUL��Jv(K�V��W��_�ړ8���/����,DU�m#j[7�B$��!�`�(i3��Q]� _�rs�i��s�٭���lC��U�T�\ ��i3�|)sՀ�T:���V�S⏸[��!�`�(i3���+�J���q���U��@����gG��ݿ�[�7C7�T���E�Ef����n`5�fK�\w��0]b!��u��X�`�ƶ��a#�f!�`�(i3�d�٣���N N�S���DP֞ /�B���a�}��ɣ�E����FZ鎬�������(���Jם����"X��[��Q[R�7E�!Up-i��e������/��$ʖT"�,�>E���]�!����w�Հ��s��&�},fcXy��q;7�B$��зq8�Ј'���Xw���,D|�|��f3��X���&RWql����g���cό���.�}�
�?�\���>��)�����_~�:N�7s�9���o>��l%i�-E�!Up-i��e�����[BC˜}1"�,�>E���]�!����w�Հ�[�=�5x�<o�;)�y��E�`JcUзq8�Ј'���Xw�j�7�������[��CC�L;Л��|#9���b!��u��c�r%�{q^:�!�`�(i3�d�٣��c�A�L'���W	ܷ�4D�P��dq�8���/����,DU�m#j[��NۥUn�Wql����g���c�rs�i�76b�*ҒT"h�p����t%��zxa(􆿳���2����.)}���/��F�z�>�/�1T[Fv�E����FWS���
�@����gG�m�D4>uF=z�{���'���>���'hZ��k��9z)}���/�}��w�I2F|:�9|X�E����FWS���
�@����gG�����욬!'B�}<����V����n`5�fK��0z�cUL���.�1�3�8���/����,D֞�Y���9��t`��_~�:N���Q]� _ό���.�1H��˧� ��)(���4s1�p#>��3���aF<��[��CCQ17�b�����$1&O^	QW�Q!r�����g �Xz���k�������۳a'[��%�э��8�>�}�����;q��b+}y[T�=qއ*|�ވQ�:�!�`�(i3K�VSƅ��	^���y���ԵU{x�j؀O��u�>����q5��'x#%��v��^	QW�Q!r�{F��#�����R.P}kBn"xz�2�w�����-����/⃓a���8�#���nh���I����{S'��⃓a���80�iN�
_�h���I����{S'���%t̓�@���{
Bk	䶙%U'��FRMv#�er�T�.@9m����1�� y��,'{w#/ B!�`�(i3!�`�(i37�wtMM��Ɇ�5�"hp��Bvw���`��״$(�>g�w�R���ykb>���p�߬�F�<��r��;i�:`�+P��l=���b��+N���ˇM|�"D5�O�%E#P�;����<�N�'t�c��B��1�^�o�\9|2I��jsz���AZ���d���!i"(<K�'P�T:���V��X�G[�q��T��|����5��"u��������f�՜�T�\ �����0[յ[+8�/w1z��ӊo�*H��&>3d?���2��HO���u�#�$IX���c�4e��_
�u�'�:����:�T�ԁ1�d �	ܷ�4D�Pt�
,c$���ޠ���!�`�(i3!�`�(i3!�`�(i3�_��U&���8��Ս9�y�ł?V�fc$��b��X���&R�n��Zn���EU.�(���[0RCm���Ӱ�e�����U|�W��eg?��v9���r����!�`�(i3!�`�(i3S`�@�t�{#	�x�u�#�$IX�b �gB�AԢ�a\�w�+ʝ��0�X:�r[3Y��P4�:5A��p��^(C<˭c����[�Y�#Q���)Ύ����X�G[�
�HYF�@��k��M�!�`�(i3!�`�(i3!�`�(i3��c$�6�byBH�}�x�gVdxQ,�,��7-oZt㧆�!F�R��X%�;���֜���áh`:,��� �e�d����\������6Bj�!�`�(i3!�`�(i3$ʩ�})�Ye�?���w�R���y�U��\JD
��_��\����
O��K�8��>L�ul|����k�5l����w����w>��Y��d���!i"(<K�'P�T:���V��X�G[�q��T�ٮ|�,
����y�<KX�+�#�W�ģI����eI�g��U-�e�,���6+���èVuD�*'��>E-�N\��be�����E8�c�r%�t^sRK1сF}���V6D�N�����,w	���՞)Ǭ�Q̞��>������*$�p/��x���6Bj�!�`�(i3!�`�(i39�O��F���{S'��uD�*'�xѴ��>3d?���2��HO���u�#�$IX��ݣ_-�1���~!�`�(i3!�`�(i3]q>�A�	����0`i�:`�+P�ސ����U��)���Y;e�iK-pm!9�>Q'݀�=��`���φ��<�6�i�:`�+PD�r�c��!�`�(i3�'ž1�|��P�:k& ��-����!�`�(i3�c�r%�Q"���_�K7͍��|��W&":�ݚ�Н�*qA����6\�4�@�� �-j�1tSjv�����l��	ͰZ����b�m��H�u�q�4\v��KVט$��}�S��J�,�����B-��!�`�(i3q�\E��0�X�G[�E�g�������(ӈ��W�!x����c�r%��S��`G��ݚ�Н��̢k���x�j؀O��w���B}�����z��>!XM�#�yP��C��?�T'����0��d�����c�r%�8�Z����p}�f������M@:��#�B� �b��!�`�(i3EOJ�uxm�ސ��� ,��rQ�ސ���6 y2��R�՝� s�#^ˤ�$����>E-�N�&Cd�c}������!�`�(i3EOJ�uxm�ސ�����nF���<�W�.�P�	��
�Q�}���%>�rGO�D mWN���%>�rGO�D mWNHN��R���IX0F�M�ꝼ�:T@�v�-�HN��R��?�d���&�af��pD���E9���T�=qއ*|�ވQ�:�t}�F��<�[xӕ�t7�L܅2�w����;����0,��3"ة�2��&����k]���/��E�u�N4��A妡��M/*�3�)�;��"q��$�������_j���m`cX�d�}�e�������{
B?�FE|���jVѭ@!�`�(i3!�`�(i3?Q�@X>#�[��N����i��T^����*�O.�Np����`yP��C��?�V�bx��yj�V��v�V\�	�=!�`�(i3!�`�(i3!�`�(i3!�`�(i3/w1z��ӊo�*H��&l���M$�[�0�7��\̍�ző�`���`f�?ǉ�=!�`�(i3!�`�(i3!�`�(i3���M$��2�w����0��5���	^���y��8=N�G&�� �(�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3�N��W��fcXy��q;d����N�fcXy��q;����pC!�`�(i3!�`�(i3!�`�(i3!�`�(i3��+g^l�>&S�XQ�����>�afcXy��q;�/m>8Φ�읣E�6�/d�G}%����3f�ZaEUԾ�� Uv@C�
]�vp�J��N0��!�x=�FZ��Q�,^-q+顳K��(*�O�q_��ҏ��ݚ�Н�t�td���5;�jmT�#i�:`�+P+鍎���a��o���H�RtV�^��l�^!Fڸ�>P��=����h�c�u��nu p��@���!�`�(i3x�j؀O��u�>����Cw�Hm�̆J�g�*~,�H�͛�!�`�(i3��+g^l���b��M�,�����b+}y[!�`�(i3��+g^l��+��\���,����"��ӌ�r!�`�(i31���~!�`�(i3x�j؀O��(�\G�@�L^�?�/��kOT!�`�(i3x�j؀O��u�>����Cw�Hm��!�>!��!�`�(i3���#�cQfcXy��q;�/m>8Φ��_2 �d���(4G��>�0]��2�O2�.+��W�Wx�Ա�%��/�qpse��\�2��s���z��_�mS8<�n�ݚ�Н���+�t2�4��A妡��M/*�3�#����R�ݚ�Н���'T���+�%�эȈ]Z����'�^�����ݚ�Н��Ra])n#���r����!�`�(i3�$�������_j���Gƻ������Ɇ�5�!�`�(i3��+g^l���b��M�-��h��ƍ2���l�!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f�`���*1ʁ���Mյ�l��d��ݚ�Н�t�td���5;�jmT�#i�:`�+P+鍎���a��o���H�RtV�^��l�^!Fڸ�>P��=����h�c�u��nu p��@���!�`�(i3x�j؀O��u�>����Cw�Hm�̆J�g�*~,�H�͛�!�`�(i3��+g^l���b��M�,�����b+}y[!�`�(i3��+g^l��+��\���,����"��ӌ�r!�`�(i31���~!�`�(i3x�j؀O��u�>����Cw�Hm��!�>!��!�`�(i3��+g^l��+��\���,�����b+}y[!�`�(i3,�˳�*C����0��G���_��b~*��s�x�j؀O��)����bX�d��-��!��EJ��7o�*H��&������}������!�`�(i3�H������"u����:/�)0�/8�fk!�`�(i3��+�t2�4��A妡��M/*�3��{��3���}Dq�f�!�`�(i31���~!�`�(i3ݑ���&�d��ҟw����f�\%�a�݌3)�!�`�(i3���%>�rGO�D mWN!�`�(i3^	QW�Q!r�����g��Mt�꾸b+}y[!�`�(i3�k��^�1�x=��oQ2)����bX�d��-��!T��6�F�",oMG~�>y�pA���(4G��>� ��A�Y�
���3ʩb��w�f�ݚ�Н�3��0���\�2��s���1�, �[���*۶&��L�H��>E-�N�&Cd�c��D�$뻜�k05����X���&R�l[�Ƶ�d�8��k�S!�`�(i3�%t̓�@���{
Be���C����/{B�!�`�(i3��F��=�?��3�����3���įէ3��}Dq�f�!�`�(i3�\�2��s�(7�Q�S^Գ3����?D�8��!�`�(i3��+g^l���b��M�,�����b+}y[!�`�(i3�����!�`�(i3ݑ���&�d��ҟw����f�\%M�m���!�`�(i3��F���K�&�a��i
�i�w״$(�>g�!�`�(i3$f��_Ub�F�S�1 �fĉ>99��j���Gp�ݓ�W���q��n-���3��Y$���F���K�&�a��i
�i�w�	����!�`�(i3l�L�`v��A�qIp��KΆ�������-����!�`�(i3�%t̓�@���{
Be���C���������ݚ�Н���F��=�?��3�����3��K�VSƅ��	^���y��}Dq�f��_��>νrj�V��vG�?-�D� ��U�_:��}Dq�f��	��x��ݚ�Н��H�����x=��oQ2)����bX�d��-��!T��6�F�",oMG~�>y�pA���(4G��>� ��A�Y�
���3ʩb��w�f�ݚ�Н�3��0���\�2��s���1�, �[���*۶&��L�H��>E-�N�&Cd�c��D�$뻜�k05����X���&R�l[�Ƶ�d�8��k�S!�`�(i3�%t̓�@���{
Be���C����/{B�!�`�(i3��F��=�?��3�����3���įէ3��}Dq�f�!�`�(i3�\�2��s�(7�Q�S^Գ3����?D�8��!�`�(i31���~!�`�(i3(@X~�H:��}�S�k�:6FY̆�<4�sg�!�`�(i3�_��>νrj�V��vN#~8"�Z�*\�x9?&�8���&�!�`�(i3x�j؀O��(�\G�@�L^�?�/��kOT!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �m�ڨ�hծ�ݓ�W����O�R�2��������;�jmT�#i�:`�+P+鍎���a��o���H�RtV�^��l�^!Fڸ�>P��=����h�c�u��nu p��@���!�`�(i3x�j؀O��u�>����Cw�Hm�̆J�g�*~,�H�͛�!�`�(i3��+g^l���b��M�,�����b+}y[!�`�(i3��+g^l��+��\���,����"��ӌ�r!�`�(i31���~!�`�(i3x�j؀O��u�>����Cw�Hm��!�>!��!�`�(i3,�˳�*C����0��G���_��b~*��s���^(C<�.�|���IkB�����X	]�k��,���^���'ƃ�3�Y1tSjv�!�`�(i3(@X~�H:��}�S�74/���@�k�F��w!�`�(i3T#�3�["���'(��Cw�Hm�̊��NM���!�`�(i3T#�3�["�7#1=��*Cw�Hm��/��kOT!�`�(i3i�Q����%�э��5)��Z^�d��-��!T��6�F���N�DNlvr5�Dѯ���-����!�`�(i3���̰�!��U`�PW}�Y������y�!�`�(i3�_��>νrj�V��v��=����%��v��!�`�(i3�_��>νrj�V��vG�?-�D%��v��!�`�(i3�	��x��ݚ�Н���+�t2�4��A妡��M/*�3�I�e���U���}Dq�f�!�`�(i3�\�2��s������x~>�"ª�����}Dq�f�!�`�(i3�\�2��s�(7�Q�#�+#��]��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3)�{6�U��(*�O�q>J�H�������>e^	QW�Q!r�����g��Mt�꾸b+}y[!�`�(i3�\�2��s�(7�Q��"ª�����}Dq�f�KK�+��o�Ƀ�?PA@?N�&�bM?��y�!�`�(i3���̰�!��U`�PW}D��ɍ��Wsp[��X��=@'ѥ���'T���+�%�э�X6و�cµ�p�ֳ�맅2�w����:��q�՝� s�#���k$ ��+�t2�4��A妡��M/*�3���X�z�q�$x=��!�`�(i3x�j؀O��u�>����Cw�Hm��!�>!��!�`�(i3�5ߧE4��!�`�(i3� ��F�����@�!�`�(i3�(R\֎u��w�`L�h��=��޵g!�%=F�=!�`�(i3��+g^l���b��M�,�����b+}y[!�`�(i3�\�2��s�(7�Q�S^Գ3����?D�8��_��>νrj�V��vN#~8"�Z��mU���p�8���&�m�ڨ�hծHN��R���
�Ŏ��Fr��j�W����H
�=�Gs]k�WM��qXt�iH��{U������0�X:�r[��J��ۍb�o��_�Rv�䩲$����#��i����+�^n=\f�5>�OS�3M��e`�!��:�r$ɓǉ�.y�U=������&G�wӨj]h�u�#�$IX���O����{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r��u?�:�H���z��l t�w�@�������&G!�`�(i3{U�����%ϨEѠ� ,��rQ�f��1.X
�:qEp�;�P�t�5fĉ>99��A0ok�׹�S�C��-<o�;)�y�5���)�ꢤ�Og<o�;)�y���:W�����t�T��?E-h���U���e�?�#	*]]�iI9�o«IX0F�M�ȏ֦�"�;�jmT�#�U���e��d9=���u��r��q�\E��09mh��nǓ<�ca�e��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�_��*��jC��6�g���7t��'�1tSjv��wӨj]h�u�#�$IX�E'���1r2ӓ�E��8��`�􉅕%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�	aF�o9mh��n�S�����	�ꢤ�Og<o�;)�yԁ/m>8Φ��"50[׵�c�r%��:؜*��d��)Ύ���S⏸[��F!��D�����k$ !�`�(i3!�`�(i3!�`�(i3Q� �_tt��`���`�{�Bͳ��;��|BF���3��2�L2���`p�~(�Mt�|�AS����t�T��?E-h���U���e��_	�Ƽ��S�J\7 ��>�:�xjzӝ���w3��׍�&�U��f���l�^!ЙMǿI?���Y� ��q�$x=����$���͜P_�_S:g�RMm�o��'����u��r��%t̓�@���f�\%���n,�d��{
BF����c����F��O�<��}�u嶫IX0F�MXz>� �!,��ف�ׂ�^�Zh$r�����P}ѭP��3���o��_�Rv�䩲$����E)e|A��`���φ��<�6��7�癆cgR������������ h�ҩ�x�j؀O��_���RQ�
��nF���<�W�.�P�	��
�Q�}�Ro�G/]%�z�-uͺ�s�η3G��Hb� h�ҩ��;�%�R��ÿ�����G��Hb� h�ҩ�T#�3�["��%���S�,�b�����zO�\l3�I����%>�rGO�D mWN��Ě���aT��3G�IX0F�M����m#p���\�'\��#�bә}��_`�tJeW{o\��6�o8:4�I���c�90Mj�dL���èVxjzӝ���w3��׍�&�U��f��_��>νrj�V��veK�	�$V�%��v�ڛ���a��҉�)e����Υ�d[g%��v�ڛ���a��҉�)e��r>�[I��:%��v��<�6�Q=�X�`�ƶ��a#�f��$�\%e!��"� +}04~B3��������h��`�����y_�mS8<�n�������%�э��5)��Z^?�4V�I|�;�Ojz����q�cp6Dq���e������/��$ʖTߧ.�go� �e�d���Y�ٔ����=�$�� �e�d��]�
�D`�R\���>��)����_(ɤ����M�3e0�g�c���i�L����;q�02�ok�nS���ވ��zNc5��;�P�t�5�׹��L<C%`�\�2��s�#�<���Ў���Z��R",oMG~�D�
K��e�G��{i���t�T��?E-h���U���e��_	�Ƽ���8|�U���e��d9=���u��r�助+g^l���b��M����{�!��"� +}04~B3��������h��`�����y_�mS8<�n�������%�эȏ�ʳ�(������<��b��M+�dr�������F��O�\E�W��4b!2�͞nOY���D`��W�.��A$�P��O�@יߌ��omq��.��|ȃ����qD��=a�^7�1tSjv�T#�3�["�7#1=��*�#QSU:��8���[{/;tiND�S���/9�=eSe.��a��o���H�RtV�^�\�2��s�U�)3�B6����Z��R7#1=��*����W���Ě���aT��3G4����NL���������gT�[�NN��K�&�a�0�����\�2��s��f%����x�j؀O��`������x��@��ئ�����l��U	�`�o��_�Rv�䩲$����E)e|A�յ[+8��r$ɓǉ�.y�U=������&G��F��=�?��3��)ʁ�]V!�>!���k��^�1Aj��t�35L��$
8��2�ֈe1tSjv�T#�3�["�Yr/r������
	��j�V��vN#~8"�Z����zNc5��;�P�t�5�׹��>�����#}�{�UA�o�cx-���P���Kn��=�$�Эs��$�Z;��|BkCD��9'P�:4�P���R9��φ��<�6�@a� ����C�'�ąC>��Ӛ��S�J\7��ZavP�:4�P�!{1�~���H����R������������ h�ҩ�T#�3�["����:�ͅR]<�YK7͍��|��W&":�;b�-�2�tiND�S���/9�=eSe.��a��o���H�RtV�^�_��*��jC��6�g���'����u��r��_��>νrj�V��v�f0� � ,��rQ��NۥUn�Wql�����"����YHN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ�$,&~��]�2+r�e?㙚7u6j�"HsC{΢}"�uf�W��Y�.;�ܞ\�x��OG_�x�S�ӄz4�m�\cw�Ϊ�z7�Qu�	�'T8�	��N�����?�d���&���V9{)�%��%��ݛlI��m�dN�<@Iv��nt=:���/z*x�n;��|B��q�gk�Nw�?��3"�9�3��n�b����4��L�O]'\gWg��	�Z�kfcj��r���iI9�o«IX0F�M�ȏ֦�"�\���F�`y������T�8k��.ͥ�H�RtV�^�}��u@:E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv�yo���_$���U4����#=��-�����2��}��3�|* ����&�*楉��%>�rGO�D mWN��Ě���aT��3G�IX0F�M�}��u@:\�	�Z��}��u@:s��� �IX0F�MV�ҁGG�K�BN
\����+�^n=\f�5>�OS�3M��y��>>�����qD��=a�^7�1tSjv�EOJ�uxm�7u�T�M#dK7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK��|<��r�*q9���%�a��o���H�RtV�^���s�`��B��cf�`7�X��=�$f��_Ub��7��G_���;�P�t�5�׹�S�C��-ְ�WA��'g��В&+��[N3Y��P4v{��lw	��m�kb㳒-??��$ō�Zm\ާ�����ݚ�Н�!�`�(i3!�`�(i3�}��u@:'@a�*�fcXy��q;�/m>8Φ��"50[׵�,��7-ZH��s����)Ύ���byBH�}�xާ�����ݚ�Н�!�`�(i3!�`�(i3����a��҉�)e�����꓅A!�`�(i3!�`�(i3P������F�zḁ�f�\%�e�
?����X���&R�ǎ)�2fcXy��q;��7<�?҄\�2��s���1�, �@F�o�6:�Γ�%:��n��D�,�H�5&D�ˎ�IX0F�M��h{���kzY
�g,\\���>��XKH��Κ�p�H#�#�>&S�XQ�W�}�.�]!�`�(i3!�`�(i3!�`�(i3!�`�(i3w� �O[s���?8�F��p�H#�#��^���;�2�d�����6��F!�`�(i3!�`�(i3!�`�(i3!�`�(i3(@X~�H:��1�, �%I�O�W^ЙMǿI?q��!��\!�`�(i3!�`�(i3!�`�(i3!�`�(i3�(R\֎u�=7�7K�P?$���Os�{��ҽ��"�.Y���5k��<&��èV5�v��cg���%�#�"_���ޡ�K���b��r˾����^n!�`�(i3!�`�(i3
��axf/����Z�S����p��~L��l�^!ЙMǿI?��6�a��)P<�ܓ�Y�wӨj]h���z��l >c��?�̒0�.��Y���y��lD�u(�v���X�c�(�M�!�`�(i3��;��L�ז�1�, �g�f�p~(ŐV(MH��C��|���8!�|!��[��-����!�`�(i3|��sQ�G����7E�׵��vH<�6�Q=��[K�9MY�^�9�Δ
w!�`�(i31���~�wӨj]h���z��l �"�Mg�ƍ2���l�HN��R��bP�63Z�tq�\E��0T����q9+t�}/�"����8�Ϗ+�8l�″*�NZ!�`�(i3!�`�(i3	�����H`��Prm!�g�x^ȓ�	d�ዪ���l��	ͰZ���H�\�{\��ɓ��wk��cN�0ׇӭ�ѹ�+�t2��iK�D�b=G�6�!~�̒0�.��Y�^ͣГ��
�:qEp��E�7e#�!�`�(i3(@X~�H:����dܟz�-��h�����dDYrW!�`�(i3��Ě�����}Dq�f��%t̓�@��܋�n焞 ����7�8#һ�����ű�8� ����iEV	5n�!s
9��
�c5ew�|�;�Ojz���)e���d��-��!M�2*详p*�з=V�Q�� h�ҩ�?V��j�cC��6�g��3�J��~mM��%�p@�Y(��<���0��´�CN-�*o"���X�+�Ra])n#���r����q�\E��0�p[nۈ�q9+t�}�ݚ�Н����F��O��ݚ�Н�;�j�����ۥ�Y�mn�	u�!�M���Tf���S�0����;�
Ҷ�a�6�B��A��8�� ��������SM0.�q�\E��0T����q9+t�}/�"�����dZG%X�″*�NZ!�`�(i3!�`�(i3	������R��CU���/ p4ZH���+�̳�Aڬ&W��%�э��XW�G�<a��o���H�RtV�^q�\E��0ÿ�����n��뾦�!�`�(i31���~�wӨj]h���z��l i1.��2����|e"$f��_Ub�F�S�1 �i|�rBY�",oMG~�Յ$�O&�#o�]�ʄ�< �SS@�
�رjwc�';��#j�ݚ�Н�EOJ�uxm�}�Z��y�&TL�b��!�`�(i36S� �*���8�� ��V���ޕe`�!��:�H�����\�2��s���1�, �y�`��vN*���k� ��$J�L�l:�
d������&G!�`�(i3(@X~�H:����dܟz�-��h��ƍ2���l�՝� s�#���k$ ��+�t2��iK�D�b=G�6�!~�n��뾦�!�`�(i3��Ě�����}Dq�f������!�`�(i3;�j���и�@�f����$�\%e��}Dq�f����̰�!�Xy|�WCw�Hm��/��kOTfĉ>99��A0ok��?V��j�cC��6�g���8���$��}Dq�f�Uj��KN��f�̰\�!�`�(i3!�`�(i3��LD��C��5��R��~\C�~��/�ݚ�Н�@v��e�ȉ�$J�L�l:�
d������&G!�`�(i3��Ψ^>S �e�d��������ZAL�:�t��q�0e�#ua9�Ϙ8�v�����(�Ǔ�`��;�!�`�(i3u?�:�H���8��Ս�2V] ,TQu��r��.Y΄�l�j�%t̓�@��܋�n焞X��ͷ(�-���|e"���Z߃2;�j����E�
 þ�b+}y[!�`�(i3q�\E��0T����q9+t�}�ݚ�Н�WH��E��E���r����!�`�(i3�K�&�a������kO�q9+t�}�ݚ�Н��wӨj]h���z��l 2�����4ƍ2���l�!�`�(i3͒t�]��/",oMG~�Յ$�O&�#o�]�ʄ�< �SS@�
�رjwcgWaU �IH�RtV�^!�`�(i3��M2χ����a�״$(�>g�!�`�(i3�Ra])n#���r����!�`�(i3��M2χ����a�)P<�ܓ�Y!�`�(i3fĉ>99��A0ok��!�`�(i3���F��O��ݚ�Н�m�ڨ�hծ!�`�(i3�n�0�I](�,�˒�;j������2�H�
!�`�(i3�(R\֎u�=7�7K�P�"ª�����}Dq�f��2��}�����U!�R�-�_���|e"����l��
*kB��`x��1�, �g�f�p~(ŐV(MH��C��|���8!�|!��[�B� �b��!�`�(i3?V��j�cC��6�g��3�J��~m��}Dq�f�՝� s�#���k$ !�`�(i3;�j����E�
 þ�b+}y[!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�t�2��}�����U�=�⳿P��}Dq�f������!�`�(i3�(R\֎u�=7�7K�P#�+#��]��}Dq�f��u{*�C<��e�����(�G�$�)�a��o���ԫ[=�.n��wӨj]h���z��l 2�����4ƍ2���l�՝� s�#���k$ �H��������0��G��e�������5��X���+���b�6��R������� h�ҩ��wӨj]h���z��l 2�����4�?D�8��՝� s�#���k$ �wӨj]h���z��l 2�����4ƍ2���lĉ��%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3��M2ϖ�YX'�(=)P<�ܓ�Y!�`�(i3;�j����E�
 þ�b+}y[���%>�rGO�D mWNG�&ց�*�&��j���3��Y$�(@X~�H:����dܟz�-��h��ƍ2���l�q�\E��0ÿ������I����~u/��kOT?V��j�cC��6�g��Wç��H@<��b+}y[�2��}�����UF��)P<�ܓ�Y����1��ݘ����$�)�vx�?.8h�.�<�..�4����Y<�!U��� '+�V�6�J�J���;�Ӏ�D�ʵ�b���n>���+H���v��έ����u���/�(�l9n�Swx�x�K_����D�;�	-
^鰺e�����U|�W�˻{Zٜ=bff{�k�(Fj�V��v�Gj7�uz7���e%�v!�`�(i3!�`�(i3}Y;�jn�R
�u���@��~h&����(Aw�,��~��A���A3�p��(�g���S�
��R/�fcXy��q;If�b����|YOF@�*���k� ��$J�L�l:�
d�P}4q����!�`�(i3?Q�@X>#�`�4�ԛD�\!����JeW{o\��6�o8:4�I���c�90Mj�dL���èVxjzӝ���w3��׍�&�U��f����vo��6�^�!�`�(i3%��v�ڹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%�������&G�H�����x=��oQ2w���B}�����z��>!XM�#�yP��C��?�LO��??\�c)���)�G��\���)e�����R�\w
��R/�fcXy��q;If�b��>!XM�#�����0��G���o=�>
̹���[�ɝ��ϳ��ٜ�]A����2�2��8��Ս��Jk����;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�2�����]�2+rH {��u��]'\gWg��	�Z�kfcj��r���(&�L��'ž1�|��P�:k& ��-�������̰�!�Xy|�WS��Wc)P<�ܓ�Y[յ� \s�{��ҽ�!�`�(i3%��v�ڹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%�������&Gݑ���&�d�����l���}ϴ��ۢ	:j�����dܟz+�dr����i|�rBY�ЙMǿI?��g�F��60��d����|��sQ�GGE�"R�ɭ}L�����U�����%�1tSjv�[յ� \s�{��ҽ�'�^�����;b�-�2�n�l3D�.������l4N�J�ף������&G��6��C��|���(�����!8#һ��ز��y��lD����HF�3ח�ͣ��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�Y;�e�O�!�Xy|�W��o���t��]�'��e�s�ЙMǿI?��t?�@�Y;�e�O�!�Xy|�WS1�ӿ�Q�ЙMǿI?!����a�}c�n��`��X���&R�B���2Lڥ����ȾmyC�0kc��g���Qrf�Va�ir��_~s�8	0X��f*��<<��lpЙMǿI?��g�F��6JJ ��iG!�`�(i3!�`�(i3���[�Q����U4����#=�Q��s�s�{��ҽ��d��-��!��KVט$����dܟz�L�[\�"��X� 2!�`�(i3!�`�(i3���>���}�Z��y#o�]�ʄ�< �SS@�
�رjwc�gVdxQ,�K�&�a�/�dI{�W��j�[O����k$ !�`�(i3!�`�(i3G!���e�w���ZxHk��k�z\b~*��s�02�ok�+�g��{��6k_ۥ���e�����U|�W����f��!�`�(i3!�`�(i3!�`�(i3�F���ᘮz��l t�w�@�Ԁ����2|Q�-l�;��5��t�;��Cٯu�Xy|�W0/0`9N1������g�`:,��� �e�d��?�1�S({.!�`�(i3!�`�(i3!�`�(i3��+�t2�4��A妡��M/*�3�ܬ��H`�쮾�\�i\!�`�(i3!�`�(i3�N��W��fcXy��q;���nD'���e�����[BC˜}1�h��N�M��e
� <"w���Uŗ�4�=+�Q��s�s�{��ҽ�1F#�֞q��KVט$����dܟz�X�R&cE���X� 2!�`�(i3!�`�(i3[:���[}T����d��-��!M�2*详p*�з=b~*��s��(R\֎u�{��b�b�*�eu�j�~ q��j�J^!�`�(i3!�`�(i3��yb�	��q9���%�b~*��s�!*Ĭ�����|�x@�iK�D�b=`u0�F��a�\#���Ƹb �����(R\֎u�f}���� �p��%!�`�(i3!�`�(i3��ӷ�*[D8�82�oFC��6�g���d��-��!D���{X(���[0R!F�R�|��sQ�G����)�
��V(MH��C��|���j�֎��](g���������l4N�J�ף��H�2^�/3!�`�(i3!�`�(i3��+p��qR��e�����P�Bmܶ��+g^l�>&S�XQ�EM?�ۄ�G!���e��dZ��@O",oMG~�>y�pA����v[v%��%�э��XW�G�<b~*��s��嶬=���X���&Rq�A��Д��u��m�byBH�}�x&���Z����h{���k�XKH��Κ1F#�֞qD���{X(���[0R\�7��v�(R\֎u��w�`L��5�W��L�o֜���ݚ�Н�!�`�(i3!�`�(i3��ZhY�N��-fcXy��q;t�;!��Q�km�������.���_��eAV��2���H��X���&R�\���8fLvރ�d�,����I{�\k��Q�'r��9��t`�W ���t�1���~!�`�(i3!�`�(i3�_��>νrj�V��v
���=b�w�����ޤ[QG�