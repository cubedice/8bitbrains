��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω������?9|[�,HJ
Κ�P/�u�x�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R��
�n�T�+F��W��`��;�É_g�?�H�.J"����U���T���딣0&_���X0���2|	p��rw@	@us���)�]&��_	��u|��yq�`݊�|���"rG�
���}�\�bJ(9�{��r�H�����طǪh��p��U>?���>�`\��Yi���u����l�|���j@��"�O��$� ���xI+r�� 0�D�A�f�mXׂ�(ѳsv�`�S��Y�ix�P�Ra����+��a̞w���{ֱ@�W�8d4؇��2O��'HY-���m���.GJ����1o���Nx� ���������	x]�<���e��8�t�~��,�O�W��s�!5�S��H���)��������ҥ{E�?HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"��-h|,���(����>S��ә�����/�4�}n'���a*�x���� ����ޙB!7����ˉ�1�:�Ω�>���h���|&���ukh�ª9���$1mt�iZ]XF��������;-;*�7��RTW�������&��J�1�KB|1<\w¹��<d�k�c��`��Z�>)��p40�zɈT^�`T�W�88�;矷A( ����_�h3��{I�B�+�7m_T���Q��K�����JU<o^.K�}G��k���؍��R��j�.(Wx*|�\m���@��O���Z鎬�������(���P����ˮ��lC��U�T�\ ��oR��m�j�.Z�wa�ҋX������S8�J�]=��R�^Ƒ����"X��[�d�a�4$�[�л���7v�ј�"��Z鎬�������(���`$�P.eE���lC��U�T�\ ���A������ml̮�7G#+�Ǘ0z�cULjaGkƊ~F˯�+)�"j���b7|#9���{k�h�+��q)F��Z鎬�������(���`$�P.eE���lC��U�T�\ ��+�_0c �w�)��O�ҋX����>��l%i�-�M�g������{l�f|�ό���.���|��p��h�d �'���Xw�E�i�m}6*�3���f�]�!���D��L#�?���&g�m��+���J q.GJ����~s���^��ɀ�Om�����67�a��c���}��D���(��z�j�)�q��1�:�Ω�>���h���|&���ukh�ª9���$1m�s��d�\l</�'.�w-�G��HZ��_V�VG�88�;矷��N�����?�d���&�<��}�u�?�d���&����}��6�v'���a00��܀�������!"���	�wT�*,��[��7%^G3�ai����3a���I���;E�@R����������S���� "5�]��'T���+�A?Љ'�-{<qH�~�!�`�(i3!�`�(i36�ŏ ���.��?e��B�'��a���cg3/F�C�����F�� 0�G!�`�(i3�b[�u2�Gp��bە���B�'��a���cg3/F�C����:�,x�~!�`�(i3�b[�u2�Gp��bە���B�'��a���cg3/F�~f���|�H.z!�`�(i3�b[�u2�Gp��bە���B�'��a���cg3/F�~f��
I�Vd��!�`�(i3�b[�u2�Gp��bە������l��I�7F����x��B5�!�`�(i3!�`�(i36�ŏ ���.��?e�#2\z���&�3Z�K�!�`�(i3!�`�(i3!�`�(i3�V���37�˱�5ǣ©���<�W�.�	*}���!�`�(i3!�`�(i3-��U��p�K�{R�^Ƒ��f�?ǉ�=Z���ֳ��m�,�0��!�`�(i3!�`�(i3�X;p`�Z��u^o"�
�cc�V��ݚ�Н���b�-W��^[�΍�>!�`�(i3!�`�(i3���K�7��6ъ��L^�t�"hzf�?ǉ�=��4tBu6�]���~!�`�(i3!�`�(i3�X;p`�C��[���ԗ��6%�a���!s�;�����)�ak�m6!�`�(i3�&8�,��i��F�ef�?ǉ�=��Wʁ���p�B�E�!�`�(i3!�`�(i3�X;p`�5�8Cl8R!�`�(i3�.��Ԕ�	���ZX!�`�(i3!�`�(i3J�]�R�Ї�J}�!�`�(i3�.��Ԕ^�|n�M�!�`�(i3!�`�(i3J�]�R�Ї�J}�!�`�(i3!��I\+��M�a5��|���瀆!�`�(i3��L	�����T-��/��@������1�so��d�a���A��`�c1+����@|ZGb���5+SC�@�ݚ�Н�����o��)�ak�m6!�`�(i3!�`�(i3�AQ�0G�F�r�f�t��5Z��~�Y���(�M����H}R!�`�(i3!�`�(i3!�`�(i3B�O�%J(�
�cc�V��ݚ�Н��/+mQet!�`�(i3!�`�(i3!�`�(i3X&|a�#�I7��-5��5Z��~�Y���(��U��?D��!�`�(i3!�`�(i3!�`�(i3�F�7��Y�
�cc�V��ݚ�Н��#�@�o0�&�v�x!�`�(i3!�`�(i3/;�Ly�Af�?ǉ�=��<H��(����O��B�r��!�`�(i3�X;p`��,Wc��I����ܗ�J���� ��A?Љ'�-{<qH�~�-��<�ξ�\zdʯ��V���ҀL���Gk��,�:�N�*�xY��j3���������g�Hn7�(��B�'��a�UP��v��M몴PBoT�ݚ�Н�U�A����;Ai�7���&@�W/�s�٩��� Ī��(�����q�ށ �~�tU^4E�}:����p���hy���N[��C���*[UxG!�`�(i3�v1a{J��Xfچؗ�rs�i��r�����[J��nh�D��'T���+�iA'R�	g�%Y��̗0z�cUL��Zi+�E���s�!��2��}��g��9|P�wAA�Ɓ=<�W�.�P�`��l�\m�q�\E��0��댁HR�\cZ��2�!�`�(i3�FQ��O�ğ�%ў׫h�JZ�lG�E
b�+|�&8�,�}6��d1��ݚ�Н�|�� Cy�6j�"Hs�Cx�V��n�#�(㷾���E.t�