��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�=A���>�LZ*IV��ӓ�������]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R����h�K�5���� ��1�:�Ω�=A���>�LZ*IV��ӓ�������]��;�I�����)O��Ξ4�"�\�� ���K�O�{����a�s�O�ET?�(�c\֣�I��B���t��|U|�/֚�?d��Y�Y0V�MG��U�;�\����vg������W�aeYgA���z�Ś��
��H,7f�t�뾌��lr�)OI3��(�!����Y�f��a�Z��V���a�\�nq�M�4�Tڢ�]�
4��`DA�rS>-�v�ﳨW�M�1<5X�M�1<5X��[5:q��?q��QN���[5:q�	�
޼���G���s���d�S��U":n�Kv!�`�(i3":n�Kv!�`�(i3":n�Kv!�`�(i3���
'�Y�z�Ft�fz�Ft�fz�Ft�f�N�uD�z�Ft�f�N�uD��N�uD���Q$D�^!�`�(i3!�`�(i3j[,F��&�!�`�(i3!�`�(i3M �̦�P�ׇӭ��!�`�(i3���s�lI!�`�(i3!�`�(i3!�`�(i3������!�`�(i3!�`�(i3!�`�(i3!�`�(i3�M��Bl!�`�(i3!�`�(i3!�`�(i32�����Vcds£����&��ea�8���	�~����a��+���L|�w.j��6��H4�
� �AH���g���	r��ܤ�18��"���] ��F@�4%�����^)�r���M�˿_��h���O�`D��#�Bk�v,�ı{y�
� �AH�|D3�M�������W)����VIW	I��?G�~�MUs +������\���T��U	�1�_u���*����	�����	����LO9� �Ŭ��2Dm�x]��.] �'9�����L.��6�H�.���2/�f��=V"N�^{")8�*I�ց��6 �����Y<�zd諒~����L.��6+Q)?^R7D�y�B.h�hC���(:�J�5`xt��R�m�!=�y����h�}Jpv��ư ��/��c�Zgs=�\o?�M��;]�Xa�v�Q�W�%-C��oW9{:n���;u���7�r��b}()pxt4���J4xʆ�7���I�9���1� c��(�U����	x]̢/����w�P����>�]!�ՄN�Ӿ��)�$�����PГ��0�w&��EO�{�������E��sޜ��*�c�N!ͬ鏈wƠ��ѹ?�����qU�%��Sr�'hJ�.;��L�OT�+?3�l� c��(�U����	x]�<��O~��#?���/�[��lq+"3��
f���&}Xa���qd��.�wjX5D	1�% �DZ�k�8���҆�|n���)kd&Z0U%x�eƐm>G�I|L6�x�+ME�F@�4%��
,澶˚C�{eC�����L��xScKE#����+�^����K�^������7�j�2>�Z�kˈ��L��i��,
o��L��j���db=�,>���iE��g�cKE#��΃��ۏ]�,�DZ�u��w)�S�3k:�(�-p9�AE�M)�B���0M��=#�V$����Oh5�6�:�����`�!k������i��f뫣J"�٫On�AN�.}��8�"풠���{�;¬>P�2-i_�Zz��$��c�g�U����[$5���k��No�v�����_���MՕ��%I)��k�8���҆�|n��T�{ ��ʥ�xw{���Fe����J�Й�m��/K5r�����}����Q������k�8���҆�|n���h��C dw�J�}d��Uxn��~�>��vK�F@�4%��%dZ&��Ǯ"�lf�~��m���w>�K�6���	x]�<���e��8�t�~��,�O�W��s�!5�S��H���)��������ҥ{E�?HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ���AOge���,I\�Z˻r���V�>!�/�7��u���nEAJ_�'��P9�L�Xڈ*-}|��ι%9��oGo�Z�J��ݪ���AOge��^\��Gx1%�^�&d�A|?_W�\I���aC�h�>�N{a�9O��Yk"1/р�{:��'��F�N~Y�9���$1mt�iZ]XF�������̘�иܖ��Q�P���O ���3�ҺIÙ=�H*.�PS�������Dɵ�p�AJ�e�$�� nU�IÙ=�HF���m¡p~z�r,����� ���3�ҺIÙ=�H*.�PS���ct�:��RE��]n�� ���3�ҺIÙ=�H<z,Ҽ&�כ��p܏�<
DN��Q�^�y�zL͊�q���Vǃ����B�6�N@���k���E����F�'n�^0o4M,�����t������ݪ�򈟆�������\�vņ	N�1�.�]V�H7'�5�}�]���!�`�(i3x�]�V���	�?�ki%�7%1�e)s 3�:��)�[���6"�,�>E��4];ˍH�,t����t�i�lK�I<��fҾ��9��ЂDa��(o��0��7Y%T��BPe.��xu	�>��l%i�-�M�g����!�`�(i3v�ј�"��Z鎬����F�71�B��>c��?�"�,�>E����-��%Mό���.�q�\E��0�����?x��#��]����������ݹ�0�����иܖ��+V.���w¹��<d���lC��U�T�\ �͹g}|�H� 7�J�[&e�l�����-��%Mm�jp=�>��o�
�v�ξ������eiy|��!k�R�^Ƒ����"X��[��Q[R�72W���R0L�>��0�]2�y�Z鎬����
C��8q��f�kN�ı���}J�|���|���O�.��_$��Y�7#�xI��W��_�ړ8���/�I<��f��tN2s���(����5���I�zI.��1��b�
~�d�9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6ea�8���	�~����a��+��uq9�����g�,P�n!K��tf��
_�n�@/%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7��ct�:��RE��W��_�ړ8���/����RY��[��Q�՝�i�(�S���N�؆�B��W+`�x�oP��@t�&�e�5
��Ib����rs�i��@�N3,(�����ϲ�CyW�f�tR�wX�ծPt�e'J��\|YX�<I@1���t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s��.|Z�����8��';�¬pX��g��U-�e,%�0g���[�=�5x�� �i�#n����Ր�z*���Be�2l��4��a��se�ξ������ei4����/��)}���/��r��H��p8�(�E{p7�j�pܔp�l
d�R�.��On��M��ҹf�f3'i3�|)sՀ�T:���V�</���/�u��g��.��U�e�7����	N^�U{xN��i>򞑻�8�1�Z���=��(hy��LLp�m~|����U�W��Op�ե[F�/�\��@��8�5x�|����1�Z���=��of�-CD֧�ǌo�9ct�:��RE��W� y�T�v��1���2���I��'��{�6�etԸ�7����|�������m	z1�Z���=���^5(9�։-�.l?e�>����c_����+�˂߮<ur�<Uee�,�Aٺ�Hۄ�2HG�T�gs �\1�Z���=�"j���b7���Øf}�
�?�?KYC'v���NE!/��Vh���*ܑe�W����n�4�{lGD�V�B��иܖ��A�.u�r���,DTc�~y��i3���w�@V�c�x���H@H�֦g�㎏qló��@d���/��=��K�R�hE!3�͸@����gG�r�I��!�`�(i34K�)s"e�>�������e���"}�`�W��f�(d0iV�6IWJE�\��[�B#���1���Q��ǺΕ������5|��>�N�B��3�>�>���%���e'6���;8=�g��U-�e���b P5b11��m$��O�&��;�L���9��Xv7�j�<���dW�ML�f���m���V��_�Ps;y>ִo������6*�G`Q>
����開���]Mݺ�A7X3�7s�9���o��S8�Q!��W�a�'�%~I��U�;�ӳ�R� V�p�rs�i�(Z6����ֱ�q������m�q�>1�Pq�@�0z�cUL�,j��=�Amx��|#9������+�^|���+mVU���������&<C���Aڬ&W���G��)3���'� ǚ�-�����d��R��YY�,���e�[=F��l��r���O>���Nn���g����g�0��oSi��oٷ;�fh����G �U�'1���w&�.��;�P�t�5��2@-�f���G��)9gUS�Z�n��[�_N9=rE'O�_��*��j?�4,qH��0��atN�s��S�+���@��v{�G`,9�H�W�nק��ןnh�sH��W. �9�����Yk��౉+�+��
��B��]��Qe_%r~�:5A��p�?�JY�)�Y`��jD4����@|����r�����R'cf���R�\<۳�B���m��h��7�p� ���:=�<�I��y�.����Pg��}Dq�f�fF�5.]���Ct=���m�ڨ�hծ��Ě�������������^��x��/z*x�n߼
�d�5�a��3��C�v�GI4�6@|��u��� Sf��ƫg�THnJHܩ+��bc�n7�}�!��g_��T�d gWVbT+踫g(�r� k�|6�8�Eo(d�J��:����5s���Z�����t�T��?E-h��$^(?��"��K��O.C��ݚ�Н����"sS<�0�zG�������&G!�`�(i3EOJ�uxm�3���w�@V�  ����'K7͍��|��W&":�ݚ�Н�ЈH����@�/�M�k��G<Y�dN�<@Iv��nt=:��:5A��p���aR�!�`�(i3�k��^�1Aj��t�35L��$
8��2�ֈe�cN�0��ž�Ć�T���7X���c�}�����l��=�O�-v�*_�mS8<�n�ݚ�Н��wӨj]h��_--���g|�m�ߕ�v{��lw	�����4�:5A��p!�`�(i3�u��g��L���ʗ�%�A�i�A�r��H�!�w(�y?!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �W?�;�끣�os�鮊R�<�t@�.�g3ZY�T5��܈��zNc5�V��	��y��=-f`Rg.�YP�׀A���`����oȺf��m<�E��?�d���&�t�{#	�x��_--���g���R�?KYC'v�����p�*��nސ��3���w�@V^�h۾�(z�k��E�2}�	76�&�;��|Bת"tg �+��5�V��Q��K�֞�`,9�H�W��<��Y�&l������8y�Ɋ����Z���0�.Q�Ћ���t�T��?E-h��$^(?��"��h��w��յ[+8����"sS<�0�zG�������&GV�Ո��Ú�'nBdN�<@Iv��nt=:��:5A��p��$���͜P_�_S:g�RMm�o��'����Tj��^�G�E�BS�+��U�,�P!6���r����܌;���'������C�ˤk!�`�(i3씁̛��p[Y���"��$;��션�~N�sȸ�"rR-��ټs�  ����'Z鎬�������(���kO��u��<��>��h�EtC�<����J�F���i���ϴ�����?�618�V�
ׇӭ�щRa])n#K�y؄@�!�`�(i3=��,���H̷_��yC��S8�\�w�4�'�)�Բc>ݣK�6<o�)�/���C�$�ߜZ�`.��53���w�@V[Z��.�~���Fz�HN��R��bP�63Z�t8��;Yv^�-w2M#-5�a�x��<��>��h�EtC�<����J�F���i���ϴ�����?�:BS��k!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��jm«Ҷ��'�e?㙚7u6j�"Hs!�pL_��P�]��x0?f��=R2� gWVbT+�,���XF:6/������,���eFz��^�̷ؠ*5�����e�`���;��|B�T���|��̬�O����B�@5�3t�(�'=8{���@2P�)�#��;�:���W+��W�1ΐ;D��G�
Rv�t~��/��=��K�_��5.�����d���!i��'T���+`��W#s�'�yq������<N߼�K�iN��VW!��' ���@�0�0c��L>�W��*(��3H��ieL�X+�' ���@�$� %7�!�`�(i3U�~�vmȋ��OY'���c���鿋�E~��k}����/]P�����+���LQ����$�����E~��k}����/����g�p�+���LQ��:5A��pw�R���y��[�ڰ��7f�ڭě�m������G�
Rv�@/�uw)"/��=��K�R��K<_8 _��s�֙7�}�!��!q��V���<	s/S�����g��+˘\5���jmY�wΦs� ��6��.��L�la�F�wF�,'�*;���#�b��{�.�t#6��.��Lj�)6)-
FkH��۟�z��n� ���?R �����⪂!t-�u	D�&F�WAM�Q��\@
����G3҇
fĉ>99��;��|BbeT�gC<�f���Ն"|ʼT7sgO .��0w����u���ei�j���s��d���!i��'T���+`��W#s�'�yq������<N߼�K�iN��VW!��' ���@�0�0c��L>�W��*(��3H��ieL�X+�' ���@�$� %7�!�`�(i3U�~�vmȋ��OY'�E�g�������(ӈ���m�r����I��)���W�w��fDC����^\���b����	�.8����-��1�&l����$�<�F�q;��|B���r��������o�a��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ��:5A��p!q��V���<	s/����AIe��0�U+�qbp@����%>�rG6j�"Hs��%�Zy_HN��R��?�d���&�ϪE�smy~�K���@�^����+���@/�p~z�r,]�H��掎��d���!iSd��Pt,��j�VD"�7�,��n6�o8:4�I���c�90B3v�A��d�G}%����3f� ��ߗsI���i����wFlE� ��\���F�`yx�>�+X�M?��y�!�`�(i3����o�a��L��Z�|n��>�my$�N��o�/���;!�`�(i3��hY-N�g3�)��b_X�XV�b�z'hۉ)��d�7�q�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�s�Yls��8��GM��-����!�`�(i3{��]��C�.��r
���иܖ����g���u��r��!�`�(i3����o�a��L��Z�|q����`U�[�l��a+Ĳ
�),������8��+���LQ����$�����E~��k}����/��&%�:z�+���LQ��:5A��p!�`�(i3��hY-N�g3�)��c�{I���,'�*;���#�b�>{Z����6��.��L�la�F�wF�,'�*;���#�b��O)�kv�6��.��Lj�)6)-
!�`�(i3>��iC���wP�>Q��ǺΕod'ٙ� �~��<e�3�ݚ�Н���'T���+`��W#s�'�yq������<N߼�K�iN��VW!��' ���@�0�0c��L>�W��*(��3H��ieL�X+�' ���@�$� %7�!�`�(i3Zt%��m&<�P8��PS~B;�T��Q׭n�L���/=9��9����C.�L:,��i���A��ݚ�Н��Ra])n#�������>vD���&l����$�<�F�q��-����!�`�(i3FkH��۟�z��n�*�&�v������⪂!t-�u	D�&��9o�d�E�"�m���rwӷ9J�E[�l��a+Ĳ
�),�#�T��6�"�m���r!|�α+!�`�(i3!q��V���<	s/����AIe��0�U+�qbp@�!�`�(i3�	��x��ݚ�Н���'T���+`��W#s�'�yq������<N߼�K�iN��VW!��' ���@�$� %7�!�`�(i3Zt%��m&<�P8��PS~B;�T�dN�<@Iv��nt=:��:5A��p
�:qEp�;�P�t�5!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2�$�)�vx%�уZw3���ҕqR�<�t@����,�ǰ�L}��tO��*�O�{��؉j����[�O6�o8:4�I���c�90�Ǘa��xO.C��WHe�Q\���F�`yx�>�+X�M?��y�!�`�(i34��|�]�Tif���GK7͍��|��W&":�;b�-�2�tiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3e<�Ia��la��o���H�RtV�^FkH��ۗg�Nri �� �X?�V��z��nԷ.#=��n��<	s/1�m+�D8fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx��.��vحwchp])6j�"Hs��zX�k����\v�\�b͐�	}�@�r�<Uee��H�ʱˡb�Ƀp�~�?�d���&��ꢤ�Og���o���T�]�!��	Ǹ�y85��t���]MY�~x����;_��8W�w��fDv����+���6�6����D5�|أͽgF"?�Q��ǺΕ�f�f3'_��s�֙R���Bk�d���H��H�2��z�b�4��Ǳ߁R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#Pq�\E��0����E�I~�*0�ŷc?KYC'v�����G eK�lݧ}�	76�&�;��|B4<d��
~�_��.��ϕ��q�"��Jl��q<uiF=�xo�R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#P�G�dE�h����E�IȪG:vmX��u��g��L�������<�^._�}�	76�&�;��|B4<d��
~�~���.�;��|B31F��~Gf��x��9�Mgw�� 
~�F�,���XF:6/������,���eFz��^�̷ؠJ��:����p�T82g��	��#�^�y�j�˗ߘ�)�I�����v�h�g��U-�e a⣃_B7�}�!��+��%�k<ꬺ��1����t��PЉ�Bk ���E�i�m}66j�"Hs)H��4)�>�|NU�jRV��	��y~��52�c6�kܜgVU�簦!N�'�y�G