��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����i�'������\ᨅh��~�a.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I��7��?'�q�Z\�R�F*}Ø���K�Z�I�?g�f���\X�<����8��U�/?��qᾪ���>�*z�w4G�� ��d�n}K-J��K��z������3�z�ω���D���+�	���lF72��{L�8br�.�/�d�������4�;(�GoAW�~.8%D.��n�P��<�w�>��S�Ś��
��H,7!!?�#�1�:�Ω��m��y�!��2Ee�Y�R2
�I.��	���
��;+$zi,��]*�8Pt�ө�l��`O��Ftl/�~8��HQ$��/z�(�^�H��y�@�Wx��gLE�z��P��] 	�p�K�I�i���^n����j�t�#wk٢ ���r:O!�`�(i3`�"��u[��6��2���k	��2�rq�\ŀ�<J�RzR^�g�EP�������!�`�(i3!�`�(i37p�J��PW?S�r�_�&�\S�d~p��M��gCu(o?C�����5	�)kJ#��t�{ڼ�`a37�Ă��>xvA�VG��1Dw>֯���,.9�}#���!�`�(i3!�`�(i3�d �^�z'�_ʱ��i�N��L��}��5E3�I,�D�y:#9�]�B�-����;���=���0)�Myիnň��h����]ߺ�`@�Ny.��d�7pp��8X�˞�DG!�`�(i3!�`�(i3p{���gM�k���lh�&ĵ�	ƹqE_���RQ�
�)T^�b�k�@����S��l��ׇӭ��!�`�(i3!�`�(i3��sƲ����e:��x����7>�����D/͘B���&,��*`O�4��.�V6���{ֱ@�,z���h���iI����p264!�`�(i3!�`�(i30tYK�yPVq�|`kK��I�+�:钾Ci5���y2�����J՝�K�y؄@�!�`�(i3!�`�(i3+���6>�2'5�sZw��Q�둩��n,��'�\�n�~��q"P�H�oe��C��c�S+d�J�Г��f�u�����!$檦!�*��Q�`��=vݖ6�F!�`�(i3!�`�(i3�s�cn0�u�A�qL��D24N<I8����\.W~C*B Ɣ��(J�f�w/�BW B]�pE(���B��|/~.)��3\�R�F*}�c}��uO0������=)�C\�?��]��;�I�Qg�@zh�S҆�|n��A�O�ϸ���q+-��e�K=�(5��_޴���΅iG��w+*��<�r�O��C��0������m�Q	��OZTv��x<܆�w�>��S^E�h/������oP����_et�rZ�?ђ��P^(����gi���$R���b�>�oa.4�����g<�R7Q߁�ܕ#؆{CM�P�,-e�]Q��s,�~TM�e�w�G3�E��])v;P���i)���zռ��+��~��'���m�!=�y����h�}Qd�А>*��4D�J1r�!o?�M��;]��,��K!�ۻ2�e�1�ΟÈ�bH\�a�����RL�a)8��Q̮�IdG�D�{����ș=I�
�w�>��S��1ﰒ�+��B-�v�
��I�{�5���l�D��s��=���Pju��w)�S��X3������e'��?��|:��0]��5w{����ր�&}Xa����1�Xhy�6�&=�D���i����	x]�<��O~����?��|:��8/Jm������Oh5"F�6x�_u�;���
r��d�;-0�\_5\�u��w)�S��X3�����0~J���;���L����/��Mx�G�F������.;�H*�^ݙ6b^�Rt����~��5��<�>e4�����5�w�yQ�u��w)�S��X3���8�W�J������;���L&+@��ڠ�D7n=�Oñ�3��f���RF�g�|�J٬Ȯ�2����	��A�A�k�8���҆�|n����5��K�O��hݜ��"���NH�Xg�����)�g���������R!�c\�1, V[���a~�d��T1X��**�SJ�й�c���R��'��z�l�w�C/��!��Hr�S@�O�{��	�Ƅ��.Sm#�yn����6����}�{,��WP=�Iw�x* [�~
� �AH�*��.��u� �(�Y�����rwjwB�y*"��ѕ�����	�������ƽ��S��y9o L�"��\�4�s���rH
>8Y�&�\�>&t"܈�E���h0�3an;�q�ma;4�2��s�D1�������v!F�_�u��w)�S �J���vy7��Mv�95�KP 4Z,^�9���	gџ�_�v%��э� �+�4W�R��Q��ȎC3	^Yt��m�ep����`�Ũ������k�8���҆�|n���f�S�z���hݜ���5��w��s�
72�5]�V���d��(3s������Me� ���Eq�iV�*$j�G�K���'�sޜ��*�D��s��.2R�Q���\�4�sW c`k��8Y�&�\��B�6��]�v�M��&�~�MUs �{<��h6���'o��*b&t�Խo�N#�_��ΙI��\�7���q���zm���u��w)�S��X3���7��Mv�9����Dtr/���zbl�џ�_�v%��X�'b�mh}����N�@N�����N���6[�'�&�' �>�u��8�F�D%� ,R�w]�y�ljrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcN���HR8�p��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�/,f$�7Q0�
8���9�X���tw:g�������!
���U��G0��#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l����2�C�b��}�@���,������0��D��L���_�L����\�Q�u|v5�*�R$������d���q����c��� �7ht��}j"�,�>E��4];ˍH�!�`�(i3MP$���p�B��F��|��v�0<๸u�Ґ�eb�3���)�[���6JHn��z��x�f7﹏T?�7G|`}���@/��(�ߜ1��E����F�'n�^0o"�,�>E��� ����{7$0~'��&\VI`,�ʺ�;[��\�v�!�`�(i3p40�zɈ�Ќ��*��4.���Xt�.U��'n�^0o"�,�>E���$�F�s+���!,�U&��/�,�#�H�1c����O}����g�a!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=@^7&ģM:�5t�W?pk� �,�� �0r��*�'yV��>���_��l���׷fh����y����vG\��o�&��v�/��k�����.����$`0�S����[LKS}?���\z-ܘ�u}����зq8�ЈR���b�>��;C@������9qj�xm�N��p��ٸ�z��������� ͢��8k��T9s*ox!�Q�W��ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3��7zgN<�|�taf��P���p�Y�Es�D��P+G2�9��?���\z-��EM���
+����r"�,�>E��4];ˍH�!�`�(i3��y�s���	L'J����Rb��Y�W,�KYeu�BY{Y����H���/�����}2M�; ?9Pjp���Ă�tTL��\�v�!�`�(i3`�U+�PAc��N�wC�����էam�XR���b�>��;C@����sђN�1�c��N�w�Q^�MY:��Ok��@����9��;C@������Jl�y0[����	��N�Ae�#�k/�z�xEQN�By3��<�]�!����M[��ǢR�����N�By3��<�]�!����M[��ǢK�h-L���H�B���5�¬����"���������5	���]���>����C���N�T?w�����5	���]���c�A�L'Qī�*pY��am��	t���o����s����Z�n��[��{_8�Y��=�}�Vݨ�,bxqX�a���C154�EY�o\��]KOӺ�
�M�����|g�Y�'���Xw�P���w��:
1���Ƭ����
L'���Xw�P���w�S=e�d^�a��|g�Y�'���Xw�P���w����p���|g�Y�'���Xw�P���w�>0�֠��|g�Y�'���Xw�j�7���I,�D�y:#9�]�B��`6�����������s���,0=]^	�&xY�J��ev�mS��0M��y��I�+��T���jB�Fg�Y씤`��p�܂aQ�"6�l�:��N��;
�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h}|��XH��9��p#�7ڜ¸<�X��/~.)��3\�R�F*}�c}��uO0������=)�C\�?��j���yU�x�3q�;�i��t�V̚z��[{{N���zL͊�q���^y�1Ɇ?He�-�cݪ�i�<z!�`�(i37�ܥ��2��3Ù��i岦�%I^sb�d"L�i3�|)sՀ��UJZ_����>bL�'��Z鎬����5e �#H��6C Uؠ1����?��c_����+��O�IC­�4���O�>�k}�r���"X��[�~��yZ鎬�������(���Jbk-����'�\�n`��!��B�T�\ ��i3�|)sՀ�T:���V��'�Kխ�Bh����YW��b'�3Aih}Nw���U�m#j[+���G���n`5�fK�\w��0]b!��u�[��l�,��@.�c��]�!����w�Հ�{.[��(��r|�����Jj���Y�{'%s�:�f~=g(���B���o��+eQ`���K��T�\ �͛ގ���]�F�ܓH�;G+�ه�ݮ{�30�����ʍ��зq8�Ј'���Xw���,D�
�eM�6��`�B7d��n`5�fK�\w��0]b!��u�7�UyR�j�=l���]�!��	Ǹ�y85�����3�|#9���b!��u�s�Uo������zL�O�]�!����w�Հ��I��JnSl{�]&"(���+�J���q���U��@����gG5m�E��P�|�Ȝ��7s�9���o>��l%i�-��s=q�SbK����D�7���`Z鎬������_�,�+���<j�B>�ܰ$p��Q]� _ό���.�}�
�?�g�T�X�!�`�(i3JHn��z��ч��,1��;���o���\)۟��ʍ8X����}_������Zs���6$�X������T��}5��xs��k��:=k���@9�������u�X3���@%�z�N}�M��C�W�~�������Z�{/J�d�,2P��GR�!˙�kgw�"��I�Ҷ�=SPn������`�7��k'�w��#҃����i3<�f�Dl��6v^�u��>������\*�滨�[��Z���I��'��\�x�����cfo <i􆣥b�ˇ�h��ʔ����d}�K�X ���C�a�}5�h�;���EWr�<�v�#j�]�!��	Ǹ�y85��g1g�y�R���CI�3�@ym⬜	�js�yO�E���%�;���EWrd���yˑ�]�!��	Ǹ�y85�ݣ2oG�M7t����`���+x�r�w�c*����Xa�R�+�t�t>
x�bG�҉��ֱ�q���]p��k��~�π� �'���Xw�j�7��fv7c����n4s1��7�癆cg���\h�\b�T��-����ʥ�nr]@A�� �	��x��|#HK��X�wS���1੡�3��/ �D�k����jw!�`�(i3<�pN= !�e��0�U���U7'՝� s�#���k$ �'�PN��dN�<@Iv�L{�Q&O7�)��.t��A\T��!�`�(i3�� л���&�W&*D�WT���%>�rGO�D mWN��h�p��L҇z:b�PXF.N��0z�cUL7k���wm����㎳5�����}Y��	}�@����U)�
xQ?M8�f2����s?�j�q]��x�4y~�4�uh�?�S���/gl���:5A��p_dW�����^���!�`�(i3U /숇�à}�(-�;S5b	��T�./��kOT��6���}U��i�U젩`#FW8�	������Mj ��}Dq�f�G�&ց�*�����Tn���}���S.�3���@�7���!�`�(i3pı��0�{�
���Z��3��w��\�Wݰ�����zo�ݓ�W���i=�M4�0 L?ஹ�%���>����x�ݚ�Н�(*�O�qR�e�ˆKۀ[}�N�`2���K����f��^�!�`�(i3�rc��a���&~e�e��E{��hNi�>��܍���|e"ʁ���Mյv��N	Ղ�I8�y\��S��z���c�w�!�`�(i3U /숇�2�D���3-�;S5b	��T�.����@����6���T��M��U젩`#FW8�	����<`�"�:��}Dq�f�G�&ց�*���%�a��Tn���}���S.�3����P��6�!�`�(i3pı��0��\rY4���l�Z��3��w��\�W���b7�P��ݓ�W���������4�0 L?ஹ�%���h9V���W�ݚ�Н�(*�O�q�\F�t��[}�N�`2���K���O8ԇ�!�`�(i3:�-���w��&~e�e��E{��h8_[��e����|e"ʁ���Mյ|�XG�^%	Ղ�I8�y\��S��z��%��Pz�!�`�(i3�Yw���Ӭ]ˍ�t'-�;S5b	��T�.�7N�S��6��V(pyL0D����B.FW8�	���y���#F��}Dq�f�?�{�X�[�g�DPp�u��A�0���򴶽!R�@�6�֐�2$%-��}�	76�&�� Ӗ�t�q�l;1�!Ԝ��c���h���E�O�����@�&_E�EYZ/��&/�>Br֯���,�l�̰��g��!�qg��^��x�=QK:2i�ȕ���Q��i7N�_�wDo�h�'�t�Z�f�}��+��\��5��,bXh��d���!iEOJ�uxm�PQ%cp��g�J��X��!���;&uL��t��B���N�gl��ܬa(􆿳�OO����˝Sz��E�4.@��0pU��}�6j�"Hs,/A�|[^O�M:R	���|�(AU4T k����ʦM~����6h�����T�ǚ�=2�L-���;@�1���C9*�¢�$�xKw�6��/B����~?H�?�����3@�4�;Ύ�@�ֱ�q�����2�w�]'�-Q?9䌎�����:i.ߋg���~�26��\\��;/���*e>�{�a�\�����fZ���o ��b�FP&P"G�wk�\���JHn��z�3���<��;���EWrQ�^���"�,�>E��4];ˍH��Oo��[*������%čr�|��B���}��yzc�?bȈ֡��u*w�A�2N��n���]%~*~��f70���N5Χ��F�,ؚ��XJbk-����'�\�n��6��	���`y���ֱ�q���z�␥&sq�?��IY%T��BP	�I]���d=��¾ȼ\���F�`y6\�4�@�� �-j�1tSjv��
�t��T&��ۥ`�M?��y�!�`�(i33���ڝn��0�|섃Va�ir[��l�,t���H[W?ð��T�ݚ�Н���=�g�żפ	�?9Pjp������PN��7�v�ԯA��bu�x��ݚ�Н��H����Jbk-����'�\�n1���R��뷅Kn�;F�Q��s,�~TM�e�w�Gr͍��Y�1E�c��>ݎ�T���r͍��Y�1� �54�T!�`�(i3�$�#{dC�(��mp���Z�{/J���#D}(��26h�W�5��|��:5A��p!�`�(i3E��\�����45��"���G��#!�`�(i3�̢k���!r}<ﷹ�Q^�MY:T1�Ɓj9��jg����ΒՎ h.\���Z�
%�A$�D0w��>�4�_���[�,�/>��a�r���m�5��ݚ�Н��0�9&،��)���4�����wb���H�1����?��&l�p�q,!!�`�(i3a3@��[/�L��O��pt��1#��
��}Dq�f�՝� s�#�K4ZRP�����9�p:}�L���)	�8VڂK�ykv!�`�(i3����&��vL n9-�N*��D�x���Q���kO��u�:�HCaIMl�i;��B��}Dq�f�!�`�(i3�JO�'��Z�UT'�vL n9-�N
�T�r�5�!�`�(i3\OW�:�ݎ�T��߶Seͪ��Y{Y����H�����1tSjv�!�`�(i3�uz�#-]iyQ���4��}�@���_rS�b�8Z�AԢ�a\蟘�26h�W�5��|��:5A��p!�`�(i3E��\�����7}#�ouߗN���g�3$�J�5'!�`�(i3HN��R��bP�63Z�t!�`�(i3%ʴ�ɒ�L��C�/�y|2I��js��'Q�:�H�RtV�^!�`�(i3{[�ב�C���#�'4v~9��c�	?�N����!�`�(i3�����!�`�(i3�H����y�A�룘8�u?��I���y��lD�\K#|�t�}���zd�Gͦ�Ũ�i�/v�ы�����!�`�(i3a3@��[/�L��O��p8�#.��#�C����!�����!�`�(i3fĉ>99��A0ok��!�`�(i3���F��O��ݚ�Н����W0�]��e|)0����n�=�H����ʒ���)0�x����VY�+��I�j� �&u��r��!�`�(i3{[�ב�C���#�'4v~9��c�	?�N����!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�M;�Ղ���C�6L����&fy��I��gs7φ��<�6�ֱ�q��r�a���B8.&�Oa��{��� �[�^[{�
��ֱ�q���GH�r@�W���3���_��Op�ե[��GAџV��$�Qu��`2|`Kr�(�'
���|���0EQ�W7��`���φ��<�6�n%���H�|{��U�=�^��#�a�Ą�ԬQ����5��t�1tSjv�d0?�s]�[�oY�ՙ��~d�[��$�-�s���o�;�E����2"f0��i�����ݹ^h	�gAkI��L�~Z?�w������b�@h�Iz�q��u��!�0�	�:]Iԫ��]�+r� :��
&T���Eb�#6�b����'�q�%bI`��}N�� :��
&T8͎g��Tu��r���D������꠼*d�m'�^�����;b�-�2�'{w#/ B�D������꠼*d�m�q9+t�}�ݚ�Н�D����pG+((�8f�A������!�`�(i3�i7N�_W\&:��;�i��t�V̚z��N�Ӛo�����Yk�����R��%4��"S�F�KD�Vr[/}>5��0�:5A��pfĉ>99��R�V�"�0�
�:qEp�;�P�t�5fĉ>99��A0ok��$�[6{�!�&X��0m_"��3��a���� 3bH2�	��x�ȓM�Me��К�CL$(�� :��
&T8͎g��Tu��r���_���`[��l�,�nz����֊��NM���.��/kjK���r�����D������꠼*d�m'�^����ȓM�Me��6��y�{``���*1$�[6{�!�&X��0m_"��3��a���� 3bH2HN��R���ء�I��߸��S�Ȍ\D�nU���:
1���ƈ$#�h�I�N�A���\�rҖ�A$�P��O�@יߌ��omq�:Fa�7������A����Y��<�b����HA�'ž1�|��P�:k& ��-�����9lD��XH S����E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv��
�t��T&��ۥ`�M?��y�!�`�(i3����,��z�
1���;#o�]�ʄ�M��,����q���f�e�x��w�����q� P�G��Hb� h�ҩ�K��ft���r|����yQ�}�\��~z���ډ��%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��jfF��v��T�#��[J&
u���/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�_f�]�o��*/�|�!����>�B$�A|'�4ER��0���Ԙ�������|,��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��xc�d�%7l# ڡ��6�o8:4ڎ�\��q��~�26��\;��B�lXm��G��*�cY�~�"���ʷ������<�������V%~YqsوiI9�o«IX0F�M�xc�d�%%1��ڒ�df�L�_dj�Ï��	�l�lM�3 ��Ǳ�_����HH��"�̙	,N��>�s�,�H��-����Z��JP���K���&��N��Ưb75���J>n�	G0��p-����`C��O9���w�w:��0�9&،��F�z�8#iY�g��Ѻ�&\VI`,"#S�K�.��5ߧE4���H����}���yb��,E�o�=2�8�u?��I!�`�(i3$K���@�!ѐXM[��? �������>�3�,Iw�)�Ć]%�L���L2��u����;	ȕ?� ̍�e�!�`�(i3f퀔�����̹�d.  m�J&�?hĪ��:����D�6S�,4��Y���$73�E�eNzL�lS��V0�"#S�K�.����L2��u��l{�]&"(� ̍�e�!�`�(i3f퀔�����̹�d.  m�J&�?hĪ��:����D�6��遇K͞���$73�E�eNzL�lS��V0�"#S�K�.����L2�s�᢯��0�Lm�<o��
̹���: -Cx䪈�*

�	�D �:���_MMDV+��PJ᢯��0�݇\��"4���]�w9"x����l���^�֪P�ꜯ}Dq�f�1��3��`�����
��A�IS��,ܓh�,�[��hg׸�� �?Ct���g[��p����y��j�ɋz�����#~胁T���AG"M:}8�?
�ǈ�MQ����ry�茴������}�	76�&��A0ok����Ě���aT��3G�IX0F�M�xc�d�%E�SR|=��Â�	�ҔD\M[�]+cDy4�$�+�;K>Ww�ǟ�bƑ���&���IX0F�MV�ҁGG�K�BN
\����+�^n=\f�5>�y_ G[[��^4�H�<���"sS<GYqcHTX�';��#j�;b�-�2�͘D5���q9+t�}����@|����^a�nu4Bޗ��jw�	���|#HK������ �'����u��r���Zj���
-�J4p'�>Sq�d��zp�s��&I/��\]� h�ҩ�-�	B(�	<L Q>=״$(�>g�
�:qEp�;�P�t�5����l�� ��5%q���f�e�x��w����֯���,mk��L���R��3����'��a��o���H�RtV�^p>��C=U����]Ծ�b+}y[���%>�rGO�D mWNfĉ>99��A0ok�����F��O�\E�W��4bmךBo�N͘D5��kK�4+�ZtgQ�9OZgY����n�b[��Z�s�Uo���,ܓh�,�F*�L��!�`�(i3!�`�(i3[��>`�lM(�s�;{�ަ.ȇ����A[g<g�!�`�(i3!�`�(i3
�:qEp'{w#/ B!�`�(i3$�$���{��{�R�S�bK����b��T@����E���z>bK���ţ��N����4�@	�u�a�ݚ�Н�!�`�(i3Ǝu1�Z����M�X���˫φ��<�6�@a� ����C�'�ąd�G}%����3f��$�uGci���{2�'ž1�|��P�:k& ��-����J>zߋ��>ַ�����ƍ2���l�����g�Z��3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l�� ��5%q���f�e�x��w����֯���,mk��L���R��3����'��a��o���H�RtV�^J>zߋ��>ַ������?D�8��HN��R��bP�63Z�t��#�a�Ą�ԬQ����5��t�	���QC�꠼*d�m�d��-��!g��J�s��03�� <I�����&G!�`�(i3�&��>��q9+t�}�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��&��>��]��E�̜�&�f������t�T��?E-h���U���e��_	�Ƽ��S�J\70C.�>��V�m^݆��xjzӝ���w3��׍�&�U��f�����C؆�AZyB�"��ӌ�r�k��^�1��dc�@c�����h��-�����s�Yls�<Ԍj��_�mS8<�n�ݚ�Н��K�,ǆ�`�íN=]b~*��s�/$�ߺ��]���޵.�ۃVa�ir���ևA�'����u��r�����C؆�AZyB�"��ӌ�r���%>�rGO�D mWN;�jmT�#��j���q���f�e�x��w����֯���,mk��L���R��3����'��I/��\]� h�ҩ��l�de�����$�a/��kOTfĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹���8�2W6�ĥ�A��6<���oA�LD!�GkǤ661��������C7@�����hH��6�3��N�߿�wW��ZN����6�o8:4�I���c�90Mj�dL�{y����i�q,?5q-�+���5wȏw�*��xjzӝ���w3��׍�&�U��f�Dw\���I\��Y�W �+��!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^L�J)���� \L�1tSjv��H�������+1�;�.��1��!*��*8M*QfY�"Z�gVdxQ,"��
������� h�ҩ΀�(���0���;	ȕ?'�^�����ݚ�Н����F��O��ݚ�Н����KL���>Ht�u�UG��Hb� h�ҩ΀�(���0���;	ȕ?�q9+t�}�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�`&c�'N�j�[�6���"����)W[�ۺ�E4�$��PGeAx�M��C�Ê&1@�-?�t�J��l{�]&"(quA0�e]'\gWg��	�Z�kfcS��KF~!��;���EWr}���yb��5������ �i7�sp>�8&���I��S�J\7������ō܈��V~�w�U�Ʀ'ž1�|��P�:k& ��-������Ϟ4
T�W��%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#��"����G��Hb� h�ҩ�{���v0yfb�YL��&\VI`,�i-W����� h�ҩ�!�`�(i3}���yb���}�@���_rS�b�8Z�AԢ�a\�2}$#h6������t�_��ݚ�Н������!�`�(i3�GI�\�0�c��v�B^`ٌ���M���!�`�(i3��Ě�����}Dq�f��H�������+1�;�.��1��!*��*8��!�qgy�`��vNiJ5a��A/��M���q� P�#o�]�ʄ�Xz���N�D�s�x�|c�Ό��b�3�怜gVdxQ,ӔРq
V2?�@,��V��I�N�?H�RtV�^��Ϟ4
T�W��n��뾦�!�`�(i3�5ߧE4��!�`�(i3?��LST拂WMG��a��o���H�RtV�^��Ϟ4
T�W��%��v��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�Ms�Uo���,�د$��ѩw���]�T���A���-`���&�\D��D1��n����ݢ������쒃\&��Ϻ��S����=�Uʮ�V(Y��a��R���t�T��?E-h���U���e��>�2���u�#��nt��F�z�8#�b9���:&�>��s��n4s1�U��B��-
r�	O)�A�IS���=Djw�9�xjzӝ���w3��׍�&�U��f��a�}�$�᢯��0����$�a/��kOT*qA����6\�4�@�� �-j�1tSjv��
�t��T&��ۥ`�M?��y�!�`�(i3��T����4.�ԫ�0�	A���-/a8!�`�(i3��N�T?w*��D�x���Q����.��$����zܳX��Hpt����}Dq�f������!�`�(i3��N�T?w��OZ|��������Y�I��fĉ>99��A0ok���H�����<Df��Eʨ�`N/��R��3���:
1���Ư����z���!*��*8b�3�旅Va�irbB@�7݂�F�z�8#�@�ܫ՞�� h�ҩ���೹�C�A�IS��[;\v�a���?D�8��HN��R��bP�63Z�tqt��h�bK����b��T@���_�mS8<�n�ݚ�Н�ըa��9�(�w}�W �+��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�ȌxŴ�Đt�|�Ȝ�ɸ�0�"�˲yQڥ�#�G�1a;j�7ߔ�;�&���b����~�]��FT;z�/j�h0gV�z�>�s�[�W�'0a��0�A�IS���~c��0���IX0F�MV�ҁGG�K�BN
\���$�Qu�F��&�o�WW;��'n�^0o���˟y{y����i�q,?5qxŴ�Đt�|�Ȝ��ShT������qD��=a�^7�1tSjv�ըa��9�_�o�@^W �+��!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^L�J)���� \L�1tSjv��H����,|ފ������o����T����Bu��r��H�����?�@,��V.ޟ���T��=y��������0�ܣ�¤�<T�I��"�
�:qEp'{w#/ BH�����?�@,��V��J����(�ߜ1���}Dq�f���Ě�����}Dq�f�}I�6���N�Cٺ��#o�]�ʄ��.�L��w)��
=b~*��s�)��7��Y( z�P��x<]+dȨ��J�	�H�RtV�^w-)Sz�MB~�S;������4Yz����|e"$f��_Ub�F�S�1 ���p`-�F/᢯��0��ڎC�?�M?��y�!�`�(i3Y��8>h����z��q9+t�}�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6���U�R.���p�Tu�i r�_��k��~��/6�o8:4�I���c�90Mj�dL�N}�m��{|�v�����G4aL��zL͊�q��D2<�4j��`���φ��<�6�c��:� �����"sS<GYqcHTX�';��#j��=����t�ִ���	ɩ���@|����^a�nu4Bޗ��jw�	���|#HK������ �'����u��r��{���v0yfb�YL��&\VI`,�i-W����� h�ҩ�Z��JP���K���&��N��Ưb75���J>n�	G0��p-����`C��O9�՝� s�#���k$ Z��JP���K���&�9�ڟ,AX3�T�#_�B�ݚ�Н����F��O��ݚ�Н��K�,ǆ�`�íN=]b~*��s�/$�ߺ��]���޵.��_�mS8<�n�ݚ�Н���6��/d.m��D�Q��H������-/a8!�`�(i39O�m96��\��;�,
�:qEp'{w#/ B!�`�(i3��}��"'�I��`j!�`�(i3��Ě�����}Dq�f��s�Yls͘D5���d��-��!g��J�s���n�{ .p������&G!�`�(i39O�m96��\��;�,
�:qEp�;�P�t�5
�:qEp�;�P�t�5���aR����%>�rGO�D mWN��Ě���aT��3G�IX0F�MNۂ�k��� $)�lj�iE�EYZ/�(��"Q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcm���D�'!