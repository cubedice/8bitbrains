��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�-Q3�Y�h��~�a.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I��7��9HrbkC �mD�?=j��S
������M7\F���r��C>C�݂�N$��/���	�0���'v6�o�"c����A�&�8d�v��x�۔7�D��:�b�#�Bn	����I@beB��H��>I��4��u"%�������j)j*[��HMi.��>��'��E����F�A�y]M���y�.!/�1 T�V	�tL��	�<�A�}Q�� �P�_ߠxR�	�$F5��wx0�<����O4��X��m�� N�X1јds£����&��=j��S
������M7\F���r��RL�a)8��Q̮	�̷�\�O~�	Q�fo�Ѓ��;H����U��Pa�ѭ��xق��X���&Ê�Oy.Nk�}u�"�*���k�8���҆�|n���u� �(����X�R��2WucJ�Й�m�N�
�Mڙ��*����	.\(��i��p��Fr'*u��w)�S��X3���8�W�J������c|L��o�H����m���>�o��[��MWb,�)���Z��or�O��C��0���[�	�P���I�O�%��H$YDD�ūG�\������c��uGQ(�9��7hm�!=�y����h�}jh�6g��+��� ���k�o?�M��;]�Qs`k�sǈY���K��j�r��!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc(#`��Gcp��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�/���[ ����ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l����2�C�b��}W�����%3?���kW���;��sD���L��+�Uz�QL@�t퐄(��ī�o�D2BC��5��Yk"1/���%	v3����M�磋��w.V&��B֥����(Ҝ�qc��[��M:��;6aJVlO/8֩]=$�G�p�P�q5Uf�Z��{�OF8��[[��V��I�Ūe��1�i��ʆ�In��tX�zgq����2��̪U��֜��3,ԯ���gn��Ab�%^��|��������Q��Ki��i�����8�TP��VchT}u��Q��L(\Ӧ����ǎ=�tneX N�By3��<�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+�\.�l����"B��$I��w��,c�A�L'��!�a��5�%]���a(􆿳����^���#}�{�,�k,^+a�@IE�U����S8��<�J�QM�A�;�֋`N��7�j2�ٚC�M�����T�\ ��+�_0c ۸�Aݡ�v�ј�"��Z鎬����[�Rs&�gg�~�+yp�l�����
L'���Xw�f�VHF��Q�#<4^�c��Et��q���U�ЂDa��(���8	]���-��%Mό���.��6[��u�(��6����j����w�V�"-4��h�]8+��T�����TSN��;
�'�����N<���d�k��Yu>�G Oag�qod�֓��+��T�����TS�uq9��� �*��H�q���r�x�\�F���ANʂ�g��U-�e�:`�0&l������K���AX�ι�����v[����������k�V�6IWJE�\��[�BweUQ�>$�㶢�&-���x�����49kweUQ�>$�?� Zh�RG�p�P��\�"i躒�W�p�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e,%�0g�������DzL��L96�`6�CY���<�I����"��|[p2e�����j��vrk�;}AԢ�a\��F�dHZ�F�\Ȳ�r�r%)cA�z���a�R�wX��}�
�?��#}�{�@�m�W#�J��P���\[$Q��
�̞��>���ԜF����am�Za(􆿳���2����.���;��\T�8���ᛚ�z�Ji�xZ��j�
�iB{�Z�_��㶢�&-���x�F`���G���`y����@����gG59#�X+�ez8�US�y��Fp����f���,(���B���ި����x�3�Aga(􆿳�ټ*w2�56�����bp��1�<��P"G�wk�١��	;q��^̽1��R��ӟ-���t��W2��$C�~x���yM�/7�!�&��R�wX��}�
�?����D)��q��T�ٮ|�,
���A�;�֋`N��7�j2��tvP��f��̞��>���I�Ūe�O��; XE�8���/�I����"��L��/ߖ��aHN��7s�9���o>��l%i�-�׎o�|��96��쏲��+�J���q���U��@����gG�⊞����Ѽz�,D��]�!���|>�PQ���b�$?ҲJ�*���z��ht��R����A$�P������5d�	�+�&IiI9�o«IX0F�M\Xɵ�y�����f�YuA(�c���_G��Hb�8�u?��I!�`�(i3�d���a؅q$��.��m�f.���G�?v��� �+��R����(1l�jG�J��u�v(z^8/BtqwdN�<@Iv��nt=:��:5A��p�#}�{�@�m�W#�a�E�Rq���my$�N��o�/���;���>]&��*j2⎜�_�/}	�dN�<@Iv��nt=:��:5A��p��@h G0���˃�In��>�my$�N��o�/���; �Z�a-���g%& J�a$�Y )P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�7<(�lb����y��lD�7m�T��Ʈ+ˀa��z��2�,�$XR�QܛOcOZail������&G����l��M��/,;�.��1�eI�׾,!�`�(i3��ѯ���Z.Q�NJ�zQ!�`�(i3�;�
�Ղ�7�i'�̓������x.�Knq/�r�]/2�ݚ�Н����>]&��*j2⎜�3�}�usT�8����ӯ�2�`<!�`�(i3��jVѭ@!�`�(i3xڠ�P�D1�"�����nF���<�W�.�P�	��
�Q�}���%>�rG�@�	����!�`�(i3�;�
�Ղ�7�i'�����t�Ƥ�x.�Knq/�r�]/2�ݚ�Н��H�����kv޶Gl7�|g�)���c=���r�r%)cA/�r�]/2�ݚ�Н��B�'��a�
�oz˸�1�"���s���IK^��M�Γ�vaӯ�2�`<!�`�(i3��w�w:�!�`�(i3�'��o�x�S�ӄz4�̟�1dN�<@Iv��nt=:��:5A��p
�:qEp�;�P�t�5!�`�(i3���F��O�VA�ڦ�c4�l�+�7#���X<��Ӣ�q�ӘS��H�����kv޶Gl�e���;���^b�~R��ӟ-���J��RQH�RtV�^�'��o�u:��_x���˃�Is���IK^�H<�2�/����*Q!�`�(i3�����!�`�(i3|�au�(Z�H<�2����˦G�K7͍��|��W&":�ݚ�Н�$f��_Ub����pT�;�jmT�#�#}�{�@�m�W#��O�޳!G�p�P�m������� h�ҩΪ���l��.�B�;�ez8�US�uJR^�d�8�b(��MdGN���!�`�(i3,\ͨ܉p�u-/���y����˦G�� ʋ�a*�Gx�����}Dq�f�՝� s�#���k$ !�`�(i3��@h G0���˃�I��nF���<�W�.�P�	��
�Q�}!�`�(i3�5ߧE4��!�`�(i3��Ě���ž_�FȮ� л�" I�M�~�^��i�-H��Rd!rf��OG����߿�}�������l���||�����M�Γ�va]HH� ;�x�����j
i���{a�?j�Z*j2⎜��?��X�x��s��؄濫�L��� h�ҩ��>=���#����ӎb�[xI��&�t�BHtK
�:qEp:䩒=]'!�`�(i3�5ߧE4���;b�-�2�:䩒=]'HN��R��*9x���С$�)�vx�/���(\�M�|����G%�MP3��s�~e��D�ҫx�S�ӄz4r���IbW���;��Jw��3��⒍~���c7�m^��F�ofqm����Lh�}`H<�2����}��M���V��6gzD���FZU��υ�	���#�e���A$�P�_	�Ƽ���8|"��w6�0��ɗ��zi#Y)M���Fe��-�����s�Yls�<Ԍj��_�mS8<�n!�`�(i3�ݚ�Н��lTN��I�gw�ڢ����Q����.��$��#�_wU|�1م�_ҩn;�jmT�#ܲ�ۗ�DC�5��t�1tSjv�V�Ո����oz�N۞��n�!�`�(i3�uz�#-]ix��?�S��*��}Y�P�4��F�(=�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�u�y-<˷\��1A����>:��2�vφ��<�6�@a� ���N��ȥ�n4s1�U��B��-����A�;��27R���\���F�`yx�>�+X�[�G���K!�`�(i3!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}��}��C˥�
]��J	��b+}y[vx��c6���J����%��v���'��o�u:��_x�'DV���b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h�'�ɳ��<�6�Q=��ž�Ć�T���7X���c�}�:
��x�{�\��N�Ś�-�����'��o�u:��_x��jJ�+�rs�i�E�8�w��ӭu:��_xk\��ϡ	��}Dq�f���i�:�3>x�S�ӄz4�XƤ5_�]\1%����_���j�[t�Y81hzg�����U�._�츅��u7rv��$�m��-����!�`�(i3�����AI��Uo���?D�8��HN��R��bP�63Z�t�Jo���j�؇�M.9j�֎����-����!�`�(i3���3rnD:��FV>o Ge��d
�:qEp�;�P�t�5���aR����%>�rGO�D mWN��Ě���aT��3G�IX0F�MТKH�{?\����I2o�3Ah	)ޟ-�b�+�