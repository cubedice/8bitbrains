��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�*���g S�7���I�N<��;���Z��4d��{�
��|��Ȋ)zo1���á�K���b��j.~���m��+���%	v3����M7\F���r��C>C�݂�N$��/���	�0���'v6�o�"c����A�&�8d�v��x�۔7�D��:�b�#�Bn	����I@beB��H��>I��4�G�x4m�T
d�(b��t�켻�S���c,31�-elwB(�93;2���Zߧl4���0�?�1~�x�c,��ws�E�x��Ѭ��S���;?�jN5#��G��Qp�'���G����a�����(�I�?g�f{ì(Q[n�+�Uz�QL�]��;�I�Qg�@zh�S҆�|n���:�o�E��c�U �=m}�R�<�3�J�Й�m�R$L=����P�X�;Qn�6
�D��t�b��M
<���٪�s����
��n�NQa"_|���voU
� �AH�)��H�]+��3�U��ڿ�e�)�fr�'�F@�4%��Y�d�u��R;+�����_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hl7�Fmi�E+���WY`�`��yZ鎬�����R�LM��ħƿ�9c�5(��}���SaB:���
�vG����BP�m��+���%	v3�R$��������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ��,5/�c�����<��`U���/�<"��0�0�G�߲�R~�e�?��S9K��B��)]�_��mNc`A�qJ;���K����Ǖ#5�u���7�Y��]�IS��}-��j8HQ�?%{B��0B���]���~68K�}:g��ۺ�D�h�N�ta�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>�τ�o��OW�p7�E�W�*�m����\@%�>4c�@�8^�-�k�w����]�-r��l�6��}�|<Y񈉝��s5l��o�A
��_�b��Xw�?�b�>�:��^L]�'1�w�z���vL�vO�
�rU�?���?i����k��u�� ���$����t֬s�'2�o����"	d�,�8��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
��C�<w��>w��Z�^b%6��P�愉V�҆%�t�3C���_��߼
�dX^�	9�e�J�� m�F3�v��e	ʆ�In��tw�?�b�>�ʆ�In��t���o�E�̞��>��3Y��t�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-����_c'�E�uv�8�����*�m����\@%�>4c�@�8^�-�k�w����]�-r��l�6��=?�n�Re��k".�����(�g
��(��N�ª�8�!�!�4u�y7�D�`��_��:W����S���w���_���`�?�b����d��Y���Z�!
���<z�2
2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�I]�I�rT�8ҵ��?��׾�n��iܕ����������a�"�5F:	���.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��U(a��,)��YbIBB�S��	�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���;*��Iy'�10`�Q*�/0�b�_dU\��=Sr�@
H$��jݺ�A7X3�R�!˙�kgw�"��I��R� V�pό���.�3�Y	���R���:K���a����`��J�>�A��Z2�����開����⪂!w �����R�!˙��^kb�-�V;�.�T��n��Op�ե[w�?�b�>�"���Zx(NÍ:��"0�i��$��'Μ�J��l��`-��y��7)�
�(�;S�+&0J7w� a����c�	������V1�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcz��[���Ė�^jҔ�@y$L;����Wp�
�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���v��x�۶;�u3mY��$bR�!�"�H�}�QU���B+�0���a�\�������޳t���92"�j
C?2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ��h֏���[��j��{�W0�Ҧ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��[�iu>�$LI^y���n#zX�����N�0�/<�U��=>bMM`)��5i׈�1^��W%h�zs�a��8j� �ee><��B9'���Xw՚�છ����a�"Z鎬������	c�u�%h�zs�a��8j� �e�[R*$�s�,�TMo������a�"Z鎬�����}�f���[�iu>�$o�I��8�����G��-͕��O�"�FWy���l��s1p����^ʵx",ޫ�^o��>n��rs�i���\��_���W�A#�q���U�T���u�I��U��؀N�&jl�o2C�g�kgw�"��I��R� V�pό���.��Ј�q%
�x�P^�(}	C-l��1v�>5o�,�Lu}0����dL�t+�R�+���O^i�a2G�F���������\��:��AԢ�a\�w�?�b�>޼�\�vũh\K�5~��o����"	e��2���A��߱�jٞ���N����H�xd�BA��Y�m��?H��zh��2s��\��:��AԢ�a\�w�?�b�>޼�\�vũh\K�5~��o����"�)!=H�-i�4��}}.1��ܐW�܎a�I���開���ۆ�#C�2���_�	P"G�wk��a�S.l"��<�W�C%����_�7>�����KW,&��(���開=$��X��a����xZ��j�
�a����c�4t���d&Fo����?H2]�9e����g�F�C9�����������߼
�d=�ƌ�:$+�[R*$�s�,�TMo������a�"AԢ�a\���E�-������?D������N>�4�
����7��M�&\})����͏x�e�]�c�����<�W�C%��T{_0\w7G����=ri�{�63�SzD
k�l4�08!��vp�P}��O�����d�n2s�ȃ�`��"��X�ix�AH�k[�^��_̨����2d��S�����H�
B#�ۉ���2=�l�����uq9����o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�!�hM�-�kǾ:op�n�j{	�	Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����"��y�R���(38�b�D������B��!�>��y�3əLܒ����D�i
��$�Qu�&�<��G�jݭ�F����μ<�e<�^��XzHL� ӃV5+��:��u�Y�KG�t4~?����:=�X��wB���to�����x��y�o�!�`�(i3\����Ƅ6 y2��R���Ě����E�i�m}640�RS���$
�)R�@�6�֐����o��1��Gv䷁=sN\� ���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ��	���X���ZT.A,�mI�p�\q��+��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
��C�<w��>vW4��`�������
��s�����E���%�a��s������XP��~�26��\�o�mW���5F:	����n4s1�ЂDa��(�_�R�G��=�gw�⽒��Շ9�/�|#HK��ehj�t�����U��+��-�����y��j��kQ�gE\�;��}Dq�f��5ߧE4��HN��R���מu��� �H�0��
�xe��f���v��ONH�y��j��kӄ��{;hnHN��R��bP�63Z�t�y�"�V��5M��z�o�:�Jr�;t�/_x��.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h9��)�N6X5�_0�ū,�mI�p�\q��+��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��AX���B��r���4�G��F3�v��e	ʆ�In��tw�?�b�>�ʆ�In��t��`UNP� ��b�FP&�ꡱ0p	�I]���d=��¾ȼƸv��*Qx���˟y7�%M��أͽgF"?�+æ d;�jmT�#�G|�776����U��+��-�����y��j��k�]�0�E"���%>�rGO�D mWN�u��A�0�Ή*��a��Ɇ%5������0u�\k|aT��3GHt7s����0��'2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ���t�'��N�R��kBޫKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
����`����������
%iq	�g��w�?�b�>��]�!��=���W�N}�m��{B���T�D�]�!��`��j(&�L��IRg&��`����6Q���,G�_baR�@�6�֐<b��5^,��4��3��w;��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>�ό�\4��\�:�Pa�v�r�G2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����"��y>�W��*(��h&��*)�e4(�geC�i��.�Y��]���{,џ�Ӆ�)�o�A���l�N}�m��{B���T�D�a�x��1�L�+��8���/��8&���IH�RtV�^�}[��O��؋�se�P�X���F H�RtV�^�d��R��YY�,���e�[=F��l��r���O>���Nn���g����g�0��oSi��oٷ;�fh����G �U�'1�"#S�K�.����F��O��V5+��:�Ąk��msb�d"L���uL-���N���kb�r�y��j��kj�����N��h��]�z�[�+�ߺ��W0�]��e|)0����)�xT��ԓ�p������T�\ ��QQ�{��x/����������^��x��/z*x�n>�W��*(���Ǣ������s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڵp�+���,�mI�p��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�I�Y�^L	��e><��B9�q7�F ��`�k`3�B6SR'��2N��n���?���^�O�=�ͦ�k�P-�wC2���՝�6�R�wX��d=��¾ȼƸv��*Qx�&�R���f�+��}��n�����[�ʥ�nr]�W,�9�9x�ƭ��]�ލZ6�`��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ���H�Ѝk�f�o'
�Us�6�И2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��AX��6Lz�#j���ؾz<�hjݭ�F���E���%�a���b<�d�@�$X��յ[+8ᛂ���a�"��:"\f6za�]��}{��/z*x�nJ�1�� =yaT��z��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���y�p�)�a�Қ���lW"`oG&2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDL�����v�/��xv�3���\��:��Z鎬�������(���w�?�b�>��]�!��=���W�N}�m��{B���T�D�]�!��`��j(&�L�i��ko�$�?D�8��R'cf����T�x��QU���^4��y��j��kL1���oBΒ���PW!�w(�y?�?�JY�)�֬w�J%�H���3�}@��9�ڮW���T�Ŭ�%h�zs�a��8j� �e�[R*$�s�,�TMo������a�"Z鎬����Y8�Sv�~�26��\�o�mW��Z鎬����+�E/(��^���jeۼF��m5i��"`,9�H�Wq�71�ҁ�\�$k�Xit֭�h��O��W���hN,��@�VҒm�fF�5.]�����������0u�\k|RSm�y��cyaT��z��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-����y�CC��s�]{s-@|!�x��02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a�!^�̖g_�3����DƯu&7���F�!�� <&�M#'���Xw��`UNP� ��b�FP&���P��'���Xw�8&���I���|I�D�{�:���Qu���%��,�,
((�H*�iH��[��(��Ƹv��*Qx}�������m������E�i�m}6�E`���ʥ�nr]�b�N����LE�ZN>�4�
��+EmI��1� ��5}�Y7s�9���o��S8��@糺뾃7܌:����3Eֱ�q������m�q�>1�Pq�@\w��0]���8-|�Dp��xs�S�)P<�ܓ�Y��=�g���>��8��-�Ϡ���:=
ҭ�3�����7V!���(����W0�]��x@�������a�"�_���3���B�1�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-����RȨ�x���h�R��4�a�"����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��B2�:c�Gm�]$���~����p��+��W��5��<�>��O�J�l���d�-}L��x�kk8/H�T_(Z6����g�q����h~S܄=lx�����bLVuA��h�#� ���Jp�1jN>�4�
���2��!읕�����D����q7�F �Sup�xg쬉� }���n4s1ՃV5+��:�Ąk��m%�l|���*A&-�Ri-jI�eto�t]`!�M?��y�!�`�(i3�E̳&k6 y2��R���Ě����E�i�m}6�E`���ʥ�nr]�K؞�*/*4q�I�w�o2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �#�����lއ�n��O۬�o�W`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڲ2ꧧ��*���xoϼZ'��io��w�gӨ*Y���wYDK�ո� ��M� �r�7��:'�� ��AS̭��u�Ա�n��g�n����@Ɯ:R���!�����`���e���R��>���J��ex$^�3��m �{3�jT��&�!�Ť̚��DƯu&7���F�!�_(����@҄���G��b�i0[�S�T"�IÉ gWVbT+�|�w�佌�&��/Q[��(���Zj���
������I/��\]� h�ҩζ37y����qls��7F���%>�rGO�D mWN�u��A�0���򴶽!���r}9���/z*x�n�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-����Mw��O��]p�H�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��̷p�`��2���AIq� :�����$I�'��~������Z�߼
�d�Ii]�%��E��%*q��T��h��<�q�P}��O��ꅽ52����$�Qu��ڀ�r[s�+<yA�rU���8�:�յ[+8�r�@|�T��\��;�,�i7N�_�Z9a��q����G��)ѳ��(�NT�|#HK��P�s)B�
u]9�#�I��-������.J7h�e�Y�GhuUO'攤��Ĝ�}Dq�f��5ߧE4��HN��R��Gu�"�0�R�@�6�֐}S�χp}���LE�ZKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>ht��D-�,�;����V��߼
�dUs�6�И2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��AX������k�f�yӂKm�[R*$�s�,�TMo������a�"AԢ�a\蟕�`UNP� ��b�FP&�����c��b�Bϱ�q�71�ҁ�(���+ĕ(&�L��R'cf����T�x��QU���^4��y��j��kj�����N��h��]�z]�leT�$r�t�}iCt�w#��@��S��c�ط�¶�`�RSm�y��c�.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc߃y����,�i��8�Ӧ۬�o�W`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�߼
�d=�ƌ�:$+�[R*$�s�,�TMo���S��c���`дȣ�3�п6_G!�`�(i3!�`�(i3�|a�T�X�n���X�8���/��כ���N}�m��{B���T�DP"G�wk��'�w*_t��2a� ��Q[R�7w����\���=�g���>��8��-�Ϡ���:=��1���h�-�"Fͯ���(����W0�]��x@�������a�"<b��5^,���vQ�+PR�G�tM�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �\��8Y`�=kǾ:op�۬�o�W`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�߼
�d4I�<w��Z�^�b9���M��A���va�{����PD}#��ůN}�m��{B���T�D��\�v��8&���I���8|�L�*�g�;˺��iz;H�RtV�^zr��s���1���!��"� +}���k$ 
ҭ�3�����*����$f��_Ub�G��VO���V�®zz ���-3п��&
�a�CJ�i#�)�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h��<RBfB"z�"���0)��0�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開#���1��Y��o��5�m9R&i�|�JHn��z�c�����<�W�C%���6V���~�26��\�o�mW���'n�^0oQbA��d=��¾ȼ\���F�`yQ��%�6�d����8֭�h��O��W6 y2��R��5ߧE4��ʥ�nr]�b�N��4�� ���V�s��6�����u�G�*ZkS0��N{a�9O�������D���J7"�p�?&7