��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pEe�1����J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR���b�z�>}��������M7\F���r����&$9g8�M>PFWD#�z":���ӳ��_}��0w�\��8׋�������N���?��m��+�ڔ�wV���C�Sy6ג��̹��/R$.:&R�nU���T���딣0&_���X0���2|	p��rw@	@us���)�]&��_	��u|��yq�`݊�|���"rG�
���}�\�bJ(9�{��r�H�����طǪ��Q��.:f��7Q�TT7��N8e
�9��Ax!P�����Yl1�xI+r�� 0�D�A�f�mX׆�f�������}0x��V����*PoI:�) o�N}V2n������u�tzZ�(��L~΄gO�3���d4��3F8�B[DP ����w`q�f�
 G��	�0o��B��a�%p&�_�l�����R�G�)q�j��U�T`���N+nȶ$	��Z��Wk:�RA�����\���-UفLx��}U�� B]�pE(���B��|�(����5��-��ˋV��HG��K	0#��1]���L|�w.j��6��H4�
� �AH�c��9�ʐ�Z�<uo�gJ@���7C����]L�����Gp�4*w ���lXc��bLh��^����������k��������Lw�l��5,
S=ذ{	��3yQ�|��x��;�1JO3Ã�����r���JĠT>⺾��D��ν��[9:n�*(�����v�=�v�ƀ��j�-�0�[X�b\g��F�	9r�O��C��0������]W�� �X�ћ�R_w���"-}�@������u9l����c�=��Z=�����td�u��.tƶ�.,NY�D��ν��䲃����m�!=�y����h�}��03�#9
�m�;�t�.{�<y�%oB;sѱE��9:�Nv��?+
��+md����:&ҫ>��?B6 ��Q�SK���B+��b��?KD@s�i����]m�!I�+����=�����td���M���ѵ�Th�f�4�u�|]	+��|5��R�#>��O��n �h	;U��C4���A�5=~�A��Nm�!=�y����h�}�ԧsd9��\�l#�+��M�}�nPoB;sѱE�%2�}���g�]��s/$��dPi���{0��d#�x_ߓ�8O�_��u��RL�a)��bB���\Y>;�>��#������ZK�� 9����E��N�ɷ���5x�`���UTݟ��ڄ�]�����톋%$ ������T�]�gUQ�D��1I��~�8[5�%fB�:��͒�&z���h�6:q��1��-=���zx=\~�:hm�R�lZq w�xp6I�m�!=�y����h�}��{�F����=����W��*HQ!oB;sѱE��q�eX;^hȳ�@�i��6��>cNKK���٨%�"��QSp4��Q�&���#�ޅD�8�>+
� �AH�D�f�u�tM��RwM��Լ<�A�����`�1�L������x�Q��t�y�FrM[�_�	�� w{j�$?������ݪ���`�2�/��\�4�s���"�KlAZ�o/5�
�+l3K�1�+��W.rֹY���8Zt'��A�Z�ͽ�ͬ5�?�GƤlhJ+=��.6n����%����iR���ۡ���0��5q��ʒ2�f?���KL�����.n�2�:p!z1��,FT��xM�$i��3��U�x��R�b�3�ƱfX�����D���R�%����T��j�����n�eabZm��+++�i'��Cx�"T4�^�o�M��Dn
0l����/J}�I��u)� ��RT�u��w)�SU��T�d����|Hj`&iC]�LT����f�+���9�����}���Ň���q`�b��+M�����ꖛ�Xj��W�-c8��"p�b^�m(hZa�.f�Vr�O��C��0����D)h�{NC�5�+D�:�3W��bi�DE�AjA��]��b�4V�U��}VsTq>9+�d����k*�jZM���Ym-46���RL�a)u����X�~篟|��.��b�QlD�^\�	9����E�E����}��r�;�f�x��BP�* �^�k��t#(�0��}n�*Ty=�w�e��!��]UZ�p̹)�3Lr�O��C��0��0�\[Y���.�l�q}���w�RIS���D	�.���c��v�!�K�$`��tT^�+Z�{�?m�!=�y����h�}q��[bA%)�IY߱�F�yW��жoB;sѱE϶dFc����}���P�����09MI2׬X����]��)�HE�fśp�k�8���҆�|n��6�H7�ص#w_Et��6�h�@j��U�)�l�~L?.Ǿ��Z���q��y;�j�6�A���<�����q���Z�$�"���	x]���~ВnK8���X4�cC��Ӕu�{��Ks��}S�O1��Z ���X2tgq��a�J�W_�<׽3���=|JG8a2H��b~��.d�u��w)�S��X3�� 6��.7q����
��e*��55f�+���<�"�u$rw{j�$?���Q���p2��RL�a)Y/̹��~篟|���DB���p�%Ô9����E�����:8E�f0� �L{�^�J��$z�]#V>W�I9����վ%��>m�!=�y����h�}m�#m����#:J��1�i��<boB;sѱE��q�eX;^h��0��bG��4=�]z��RL�a)�K�6J��~篟|����dִ����h<9����E�,��{�M���o����Ȋ�څ��:;xꒌ!��S�g����$>�)]�y'��BS"�9 \D�GB<xA��ظ+
� �AH���н���(�Y���m�VV}��ԏ$��c��)L�����B��;��	k|�6|����J%�hu�՗Xr��Ӧ�v�5ܗu����q��<O}%��f����>�5%q����^���#B�zH�퇟�J��O�~���RL�a)P���6z�D�~篟|��0�Z����݇+���9����E�e
aZ�Ბ��ؤ��PUbۼ��n�/5���s��fBd:����}�2O���\�4�s���㚗���BK9�H�>�����\��)��&��U�)��NT[�z�N>d�k�8���҆�|n���#_;ʎW��9�������5��U�)� G��M�Eé�H���(L�q����n3X�$�3�^���8� ���\�4�s.)s:^�e�K+8�M�A!u���u�w/�ֹY���8�L� *����w M��b� �O��>�iJ��v/^;؊�]���c�����˘y'��BS�Sҥ��|E�EYZ/��V��$�� ��D��)��F|7��#댽5��}������2�e���6���09��U�TC�|V
� �AH�|D3�M�(�Y���mzU��ͤvc+�^\L�����^�����K�d���7U�� ���﬘K��U��+�Xa�H(�˕L�q�ع	z�; ,@�� N���� e�J�Pn\�pD��ZOU&����4����\�4�sg�oXx��U�(�Y���m ��%V��~&[#a�i�L����e��
@h�=z�|8� zgZߌ��h}��OH]_�ww�~�$��	QIe�y� ے���"ڻ<Z�V�$��?�6�b�N��D�D$���1�?1�U�<R�@.l�td���b�'Be��aWGL�y��i	3��'�al��pr�O��C��0���M�<lbts� ����Cb��W%�FoB;sѱE�B��H8����U�BwT��TE���`S���Ez2j��
�රB��uogU����RL�a)'r�Ӟh� �K+8�M8xU�?M���9B-tnD�ֹY���8�R\��G�8Ğ�2��ͧ�p1�fv;�u��w)�S����w�~篟|��� }E��R���6F9����E�t��̙}�ɨVu��7���	x]�m�Je{q���~W�*���:��!u�OMp�0V�u9l�����y�+�B���w�#/lr�O��C��0���/���k�Y2������PϭoB;sѱEφ�����9l~y<�t('�0�ɹVi��ӯ�0��\�4�sR���i1�X �9W�5\;�+^����S�5��L�����=ذ{	���g��u̘:��/�~����P�N��m����/��p������Jힺ��Ľ���~��@�}+E���Q�:�f���t�FRsyѳ����nTz�h���s�.�Jl`�X��IOb\y$�����k�8���҆�|n����Շ_ Q ���F���D�|)u�}f�+���1�*����Ѷ'��*{�@k�?o�r�O��C��0��$�>��w�	3:�y��gh����oB;sѱE��d�&� k�#UE8�T�h���:�?U��9��̵�*�&om�Vu��Y�  �[�|%��R���4����q�˯�)��FB�����o���㏞ �ب*c,R�1000��v�-�2$�z�&������P���<��2]LEA84e�t��e�×�umn��b�Qɝt�L[�il�h�7QC f�V��zK���D]�M���E��	&�~��FjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~������s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcN���HR8�p��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�//?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_E$ô&y��ѬL�1m��+Y#_WӇ�s8[ZΑ� �}E+�E$ô&y�#�̔"v��ƒ)?˳ea�8����]��
��rE���ƪϤ�Yk"1/Y#_Wӆ�q�©����0�w��7���I���}����E���ƪϤ�Yk"1/Y#_Wӆ�q�©���H��JnXe�+�Uz�QL�W*g;X~09h�i�k1i�f1?�e�Bw�M�?_W�\I���A#|��[�m���w��L�����'�@���,������0�ea�8�����B}rs���{Z85۰���N�y�g�M)ԉ���S���M�&P��yv��*����W�{}�hu��K��C����W�aUE�R�D�*��O���L KF�=B�T��%�~�5�)N�i�ĺ�T"3�����'l:}��Q ��k\�\�KE���H���o���&�t.�}��L��t�q1NJj8֩]=$���GZ>.�0�[7�d|���XP���H'˯?k_��]V�H7'�R�^Ƒ���b9���j}8o{:�����Y�V�����ϲ�[7�d|���XP��Ȩ�wl��h�U����z~ﮅ���gzL͊�q���}t��C��>�~I��M�H�ɇMk�c��`��'n�^0o����SVcU�>�6>�^56�c@��v�'rYI��RhF��j��T����'n�^0o��l���8��P�ǍZ�J�����+�'T�Д��*j�B3g�����zL͊�q����ϡ������5�hbvk~�#x��܃Ae��'n�^0o<H�-��*s ����
D�ZLN�	���b9����pP�o�8֩]=$�?�R��n�~x�9̺��\�v�T?�7G|`^�R@Κ�2e�J�Pn\��J��H9��\�v����UĒn�{���e9��1WA"SӠ�|&��6����U��+�XhU��`��&�b9����4�6�t�w�n����|��T�5�d�,W�� nU�IÙ=�H��'�PD����
q<O�n����9��#�B�sYC��\�v��_�R�G/K��(�������i{±�sR�{F;�f��X��Ye�?���j�g��$P�M	�D�$��띂ii�4];ˍH��T�K"
���d�8���obzĀY�ɡH�� �YߥթD�[*s��l=�L؅��FJ���/�`�����Y��,bxqX��b��v݋N������M}Ĭ����[7�d|���XP��ȁ<ቐ��jVM�-��(����<�r�5j�'n�^0o�i�f�C�*��M��p����d0e���c���������\{J�~���.s��l=�L؅��FJ����HwL�X�+�p}f�~�ڳks��l=�L؅��FJ����HwL�XArߟьvb^:�x���;���L��GD@�F��q� Q�e��{�-���`��p�Yl�}gL�'�����D��)A�\.�
�O�}݋GD@�F��q �VL�(\��'&S�39؍��R��j�.(Wx*��|��pe���b�c��Et��q���U����?�!�`�(i3��|g�Y�'���Xw�E�i�m}6	��	Mk�rv�ј�"��Z鎬����A��:6])�/g\�H)��,vw+�ne.��xu	���S8����ٺ?��Ʃ��6��G"ڻ^!�g��U-�ee�@Rv����my$�N��o�/���;�%ؙ,{F�"�,�>E���TD��ό���.ӈ�=�$��zigzA=v)��(�
t�ژq���U��ꢤ�OgB�Y���c��|g�Y�'���Xw�j�7��ct�:��RE��W��_�ړ8���/��@����#4� }'�8�������5	���]����,�JL���r�I+rΫ�,v���٧I�^�i�����K�]2�y�Z鎬�������(����U6�bL��W��_�ړ8���/�����FZ^�u:��_x�����	Z鎬�������(���8'qG%��Y�7#�xI��W��_�ړ8���/�I<��f��tN2s���(����5��-��ˋV��HG��K	0#��1]��N��;
�'�����N<���d�k��Yu>�G Oag�qod�֓��+��T���O'�lR�ܓ>��iכ���������N�W|�.Ҩ���"��yk��Gfz!���+��+�Ę�a2M��A���va�{����PD}#��ů��èVγ��Q�%��L|�[��܇��C��>����[t,�D���K1P���n�� d���Yw���0�;�P�t�5�a�LD�u�C�MV���;�R�I͗4�L �׭t��y(���GLo���#�hW�D$2���7 E�B��.��I=�66C�&/����� <&�M#���}�|��n4s1��7�癆cg(��_�8)$���}6<6zY~G���jO���a�6�x�?8�Bg����*F�	��x������a�"�-�L�߯v��F���5ߧE4��T2����
4�L �׭t��y(�����	w������"��yv%a��!)�����f�ƳaBA�u����`��l_��~��D�AV� `A��~E��~sv��k�6O����Ҷ�=SPn������`����8-|�D����<�.�%m,d��ߴpiʮU:夼W�F
�ੁ��@|������]�9Wp��� //�q(�HN��R���ء�I���RCz��QE�7��%	�0�q����"��yz�Pr��� �v��X����?��9�Uʚ7�ܩc�r�(���JHn��z�r��]�]��eCǮ��\�v�w�?�b�>��#�ڊ<?@	�+�&I(&�L���
Ո�C�hk��Y��A�m�(����V��J���6���ǈ-��ʮU:夈
N~�k��5i^��]B�e�x4�v�w�{C��Ě���aT��3Gr_0<����K�b�-)Wi�l�U����;�� D�4o�2d�F�����a�ɒ,��N��g()��ikp���H����b9������baBA�<om���b9���M��A���t���92�,�q~�{���+}��
8��h.�A���ۖ��<��Z@Y��[�5J�<om��1��b �������a�"����'l����w�ǻ��v�8:�83�x`s6S0ʹȎ�~B�D5�O����1;[lzRY�ȝQ�~�>����<�Sm��E�̔��E�i�m}6�LFC7�5t�O���a����.��B�M��:�گ}Y-h��!��|K�{ߝs��ƒR�j�o]�����/� �UR0�}D�)x�?{��
0#`�1��JHn��z���}��-j�U
�D��JHn��z�c�������b<�d츳��S���R*��w�ǻ��v�8:1~��vA�6�6]"%n��X��+ǅ�<$M���A�,h��W��n��th�U�CLB�D5�O����1;[lzRY�ȝQ�~�>����<�Sm��E�̔��E�i�m}6�LFC7�53{@�5H��Ve����7�hύh5�e�67���L����Ҙ$7�s�U�gi�Pg`���g()��ikp���H����b9������baBA�<om���b9���M��A���va�{����U ��z�!e���im�th�U�CLB�D5�O�X��WG ���y�9�3��|?e����hbvk~�#x��s:���<om��#Â��&?��Nj�a=�X�byA{�J*�Rs�0c�툼��#���F��3�k�n׏�����M\�.$�t�s�U�gB}�J�u����;�R�I͗��ay�Ȇ^���x�k]m��Zx�.��[k�'��P�d�X�VM�����a�"�'n�^0o:���^śe�j�;��#���F�xe���vr��_.�yE.�g|&�f�B�R���>_�?"�����X~�� ��LFC7�5F�:��5W�Cq��O;�G�Z��Y�#�{U��óM�˄No�M���R���V�)s:�������.<mjR}��ƣh���%����=Y��i��M����V�܄WD�4�\��JHn��z�c�����<�W�C%�b	�4© �1x�itk��԰�/"Yն���N�PI-%��֥��ع�����������.��4�F1����|�5Cn
V~$B��~���nr�l�L�T۳�͕���y�9�3��{�"��}&]��Wu�LFC7�5J��K�R���V�)s:����xZ;a{-�K����r�t�E�ߥq���P��ʬ1H���ih}N�}h?��].�Ч���S1$� �!%��b���á2�7�?��i,��&lG#;�:E��$vi�N;=��c8?-+eN��zʛʑS��_���!+}$|~ïSup�xg쬉� }�����v�WM�v�1a|JHn��z���P��(�鏄��m�q�»Ą �N��B�)Y N��r*�1W�V�bS�-�=q�:�G�c/*��t�	��{��E}��kA���g�AmY�f�aV6�$p��9:6�5F�&� Nm�Y7 �.�AmY�f�e�Tpv�t�	��{����f��r/��5Տ�E`����?"�����2$%-��j���;��D�2�7�?��i,��&lG�i��m�P�óM�˄N�9>�N�6^`�[J�q8w5���5��0�#j�� ӫ/��m,fF�7�1Y�ΊS&v�c��Q��"��0����E�_������h�ӵeo�i� �x}1Y�ΊS&�3
�v�v-}�	mp)��y������8�i����k!�=M]iiHC��\�v�w�?�b�>޼�\�v�.��C�y/=3\H�>�B�Q��>rM�Zc�󆱼[b�I���\�v�#�1�N��>z�Vg.N�����XF���f1�0�u���A�%��fOX���0����<om���g����JHn��z��c�Bo��\�H��/Sg���My���"~6���aq���J���������������A�\>W�/Z����_]���T��\�vś��Z1`�x�y�Zglϣw����ҤJ�;
���;���EWr�_�(�X�w���vc�f70���JHn��z���P��(�麹���1[	1��r�.Gb�TG|�wx��`��Ƈ_���˱���v�B|+�{���cn��>9V��9L%��a�e�7ٝ?��;
V�;���EWr��(Q��;��b�=�j6X��z+'JHn��z���P��(��0@ٶy�i�^�Ax�v�H�J&����4��(_�<�� ��b�FP&f�%A�)!�`�(i3!�`�(i3�a�\����ο pX�謻��������
�x�w�������������� �1x�itLd�r:ha3B��*w�C&�5,���a	!33֬�lPCrM�Zc��~�/:��ǆQV���Ҥ�������|I�W����x�A/�n6�r\�H��/Sg4�y�)@��]��0�ȍ�x�>c�K����&&\�0���eYk�	�yOx(�i��/R�Ȟ3I	��.ᬵy��H *4�ڮ���Bư��9%2�8���x�Y�+���]���J*�Rs�0u����x/��'�ĮpYÕLM�(�� 	l��lB���U%�p�zꥦ���i͑��Ԣ���C��괽���5��g����;���N��-Lk���ޟy�K����t����==�x�Yu�~����J*�Rs�0u����x/�'��ޙ4!ֱk���p�˳c��sCF��[ S��x�%�/�d�"�hm�^�6/
��VLM�ǩ��8���׷y�S}m� 2�k#ʘ4��\��sپ#�J��v�8:I�}-��^R��	�ݑg()��ikp���H���ʤ4���aHUv�׿e\V��/��x�%�B���vs.�^�6/
ڌ����S�|���#q��iQ��ׇJ�	�LÆ��/�i�����܍w�S}���d����_�(�X�<�q��Dp�$�D���O�J*�Rs�0��ٴ0_ǒ�;c3Μ(4��������KܫE��gD�b���k�%\��g��\�G����3
�v�v-}�	mpҭ���^���b��v݋N������o��^EјHo��L��}�Y�PX�)��s����,�Ğ<�q�;���N�?~h��dg()��ikp���H���s��N�Z{\�H��/Sg5����GǆQV���=KmS��3D�� <(rK�� ���Q��Q7��.ᬵy�����ܞ���3
�v�v-}�	mpع��t���f~�����"��KH����t����ǅ<~!�}�Y�PX�)��s����H�r_�[=���r���e�ĵa�,�J��/R�xTGQz�a��mHw���v!�n��ˁ4bBaZ���=kif�� ����p��}��aq���g0����Xjۙ�)��s���	f%�\G���T�qb�,�����2z�R��Ȟ3I	��.ᬵy��E:@{
�Wx$G&0ɑA���
�xϥ��Nǆ��#���F��z+s)x�?{��
0#`�1��+j��Y:s�3D�� <���Db2vT۳�͕��T�1�����VC�H���X~�� �4�04�jf���w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m/��������|O�\�+�q�� 6x�@Ts��E=��T7���j5r�n0��23��-��2j5r�n0���Z7£�&�x(�i��/R���m��g���"~6���aq��yx6�n)_���fx'v�ao.\C�k��ݍ���)�{:�ˎ]":V���"^[��G�X���`6X��3
�v�v-}�	mpҭ���^���b��v݋N��������;B��XOh��M�l3B��*w�u��mo����[`�B'�&{�zYa�,�j?Q�����͵De��2Q�����ݟ���O�͛PA,q���R�*ؕ��A�\>W�/Z���N+~�{-M�O��~�O�β\�{!ˎ]":V���"^[��G�X���`6X��3
�v�v-}�	mpҭ���^���b��v݋N��������;B��XOh��M�l3B��*w��6~)?�A��[`�B'�&{�zYa�]¬')4�5��͵De��2Q�����ݟ���O�͛PA,q���R�*ؕ��A�\>W�/Z���N+~�{-M�O��~�O�β\�{!ˎ]":V���"^Be��Dc]�`6X��3
�v�v-}�	mpҭ���^���b��v݋N��������;B�鉞(Q��;��b�=�t�}�t�&�}�vo;��|O�\�+�q�� 6x�@�	�x���!��z3�:��c��%2���ʏ!	��c��*��'�/7Ii�^�Ax񣘂D-\`����y�]��b��~���"~6���aq��yx6�n)_���fx'v�ao.\C�k�Ǆ}�tu�������&{�zYa�w�X{��̳,�bC�,�����|Iq��^`J�Ύ�&
�N����A�\>W�/Z��B���[@���[��QPw��r|��߇(���м	I���������)�>��"<�q�%,��7n�!����&A��kT��4^i�u�J*�Rs�0�|�:���@�����\�H��/Sg� c�Z�q9<~�p_�X����)ͶG�q�5Սó�Ǫ��z3�:��c��%2���ʏ!����>2{�}����q�rX�]��C`e�n
V~$��&��<+'�tL���lϏ°�� ���4^i�u�J*�Rs�0]�����sk�����\�H��/Sgf����O�9<~�p_�X����)ͶG�q�5��5v؊	�\�G���nQ�rV׃_
"Y9<~�p_�X����)ͶG�q�5�D������aq���5�*��և̾\x#�d+'�tL���lϏ�l��I�K�4^i�u�J*�Rs�0]�����sk�����\�H��/Sgf����O�9<~�p_�X����)ͶG�q�5�Ӂ���zm�\�G���nQ�rV׃_
"Y9<~�p_�X����)ͶG�q�5կL�З��k�aq���P�ۑ1A�)�{:�ˎ]":V���"^�򍝟�O�<=�3���9{lq�"�$���tuR�3D�� <�1��h>��dA�Mi�{�X����)ͶG�q�5����,?n����'geWP����p�8�$��gˎ]":V���"^�19TH����˓#��͇!*��6���;���>�T�Y�^���[KxM�h�e��SV�Cagi�"XOh��M�l3B��*w�1��~��N|��|(F9%2�8��=����T�|��/�ciJ�����'geWP����p��{9LBi�^�Ax񣘂D-\`�����SVcB�R���>_�we��3��we ��g�1P�n$~��/F��"���5ߧE4��rw�&�z<a���	�r��5ߧE4�����|u�EQ73)y	�Ȟ���p�o�QM�Wf�b E���?�Y�͎�6%V�J��5����`K�c�ҩƮ���開B�m�/gV�gK��J��;=�LT�I))����A�m�(�b9���;��/ƣ��>z�Vg.N�����w<���i��ߨ(,���"5�o٥�b9���3q��=$���A���ۖ�.Q�2�>�_������M���o�G�m�?@ux�[����3���ne66�v��G���V>�R<���.{2YX�i�R�ռ�����|II���XԮ�%Ah�%4
>��XP���v�c��Q��"��0���g���a���0i���o�)-�I��'�nQ�rV��(QH�����/��1IÙ=�H��fx'v�ao.\C�k�)x�%���J*�Rs�0m�������.{2YU\��,�v��|O�\�+�q�� 6x�@1#��Z�����XP���h�5,Wl�/�O'�=��sh�ƶF�A�%��fOX^���֮���"xC��-�T(u	M^�.�/�92JHn��z���7帘��3�=r����0�i/ȇ3
�v�v-}�	mp�5�#b��Ŀ�ġ��,��%f������s��2b�9%2�8���x�Y�?A����\�v�{=J�����cP$�̄�Xjۙ�)��s����Q�^�y�N��B�)Y����ud�h �x��b�TG|�wA���^�Q�^�y�zL͊�q����sپ#�J��v�8:I�}-��^R��	�ݑg()��ikp���H���ʤ4���aHUv�׿e\V��/��x�%�B���vs.�^�6/
ڌ����S���;���V"�Y�y ��FA��m�;n��^�����4�Cf_�~z�B�6�U�D?l5�	 ������ڝ�ӡ���<K ���3�ҺIÙ=�H���ޙ���9%2�8��"ء}�6=����t����==�x�Y�����5O�%��/q|F�W�1'����
3&d�X0���b9���JI�5r{�ŵ �-�`)��\^�#�n�L�nv\�H��/Sgn��ngF�v�c��Q��"��0�jH��E.��J���6ΓU5ib�H@�A���ۖ��uEz^��r�&U������G|M����L"�9-B���H��@!�#-�[ҭ�x��`��Ƈ_���˱���v�Ր��&��`;�nQ��%>�K��JHn��z���P��(��j��ICmA�zV���!�`�(i3�E����F�_���˱���v�`4�ōuN�2�q�]�U�J�"�3ʆ�In��t�Z�	�і��ʝZ��I5�4`UV#-�[ҭ�Rw�)�� �`��YF܂d�ۤ�|��F�����y�]��˓#��͉�(Q��;��b�=��o92�t��zh+�,�l��=5;2qa���6������1�R+-h]��C��T�J���6�&]��Wu4�04�jf��=}'t<��ġ��,̓NQgk�0�y�S}m� 2�k#ʘ4��\]� ���_�hbvk~�#x�<�b��'6\�z9W�j�˳c��sCF��[ S�=¯\��/�d�"�hmB	�"�&TK��VLM��FA�k���th�U�CLf�� ���:0>����0H�����r����q'�P3�^�P�qjhbvk~�#x�Y��vS=l=����Μ(4��-Aj����;���H�ܸ��쇰��u͊Μ(4����,��T۳�͕��D����jF��b�(� �	T�����3
�v�v-}�	mp�cA�N���^����A���ۖ���M��/o��sSYqυ��ƚ�8�v�ܸ���V!_?�q�.Μ(4���؇~,��%x(�i��/R�Ȟ3I	��.ᬵy��H *4�ڮ���Bư����!h�b�TG|�w+���]���J*�Rs�0��ٴ0_�_�C.�5��4"��B�*�A���ۖ��<��Ze�C*y=�_�n�To�[w��{Q�n
V~$��$�J݃����t������@�a��#���F{\��@�����p��}��aq���=@�w��d�bș;��D�h�$�� ��yo�}�Y�PX�)��s����A���cZx�.��8wCc ,P��#��\��v�8:HjHf��x(�i��/R�(�r��])�Y�^�8�2���H��V�ß@�_�(�X�"䉾���9%2�8���x�Y��Z7£�&�\]YD�^�O�<om�����0M�C�T7���j5r�n0��:�_�B�T�;���N��6H*��l�A���ۖ!���6�,N|��|(F9%2�8����$}ům��ࡔ 4�U����ʹ�w��r|��߇(����<5��������|O�\�+�q�� 6x�@t+%x1ef�we ��g�I�����R>��o��b�����V�I�e!��nH�W�l,ѳ��=c�f������C;ub�(��n
V~$T�1�����VC�H����X�:�8�[b%Ɨ��H�*x����=��:������4�04�jf�5ߧE4����DeH�J*�Rs�0�|�:���@�����\�H��/Sgf����O�0~+�+���}����q�rX�]�En:K��$G&0ɑA���
�x����G7���
�xxܟ�,3JWh�x#�L_����	�r�@���rahZ��c��B�����y}�4N�?��y;�j��-=����`c�6��2z�R�:�F���WըjB�B[�)x�?{��J�SqVE�e�H:�I0���ԏ����[����J�Cp�������s�`�|O�\�+�q�� 6x�@�	�x���!��z3�:��c��%2���ʏ!	��c��*���DeH�J*�Rs�0�|�:���@�����\�H��/Sg� c�Z�q0~+�+���}����q�rX�]��ulC�rs�����)�m߽n�Y�P3�lWD�Ey-��OI0���ԏc�r�(����|��I�e+'�tL�"��%�D��.+;�fQ�X����)ͶG�q�5�b��YZ~w�o���*ٝ�/�K^b�;��	+��������T�s Wd2uUrG��|�S�
���N�@E�V)�jP|B�1���}܁'A~)2	�ߑ��J�*|��������2���t9�'��_�K�z��d>Q���G&o6����V)>��O˻����|IzB@k�G,<O16�,��p���#4�Te͉�Xk<�zPӹ�&�w�򪥃�n�{��l[hbvk~�#x��d2)#^&|���BY��l��=5;�D�A�'�G�}�vo;��|O�\�+�q�� 6x�@�	�x���!��z3�:��c��%2���ʏ!	��c��*�\�G����3
�v�v-}�	mpҭ���^���b��v݋N��������;B����z3�:��c��%)���;�🏡��������Q����N�����,eS=�oAg{Y#0����l��=5;ʎ��_��I	�Ȟ�����hLKW�@u��q�q���3B��*w�N����P�}c���x��z��d>Q���G&o6_��'��堼���*��P3�lWD�q�5�=ڭ��"xC��-�T(u	M^ �(팵������,�\F܂d�ۤ�|��F��ms3M��o(ͻ� ���7���ì\��2l��͘r�qU� e��kSA\g()��ikp���H������b,Il�I))����A�m�(jXx��pM�֬�lPCrM�Zc���߀1��5�e'h�&� �th�U�CLf�� �Q�@&�?�֬�lPCrM�Zc�������֯���v�8:�tV����/��n(��N�����,eS=�oA������w2}�<��bd?�&�������]�cn��>��[KxM�h�e��SV�Cagi�"��(Q��;��b�=�U3{����B|�S�
���N�@E�V)�jP|B�1Թ��q��T\�w��V�)x�?{��J�SqVEF����#HI0���ԏ����[����=�5��@��H��@!�#-�[ҭ���Ѝ߸m��c���nJ�	�LÆ��/�i����zYק�̒�H��@!�#-�[ҭ�h�s
>5�hbvk~�#x~|���@�ճ�%)�r0z�1[FQ������-Kff���e�F�N�@E�V)�jP|B�1��-XD���FA��mӡ���<K�3*��hbvk~�#x��Ύӌw��i2n_����9��b>��X����)ͶG�q�5�ms3M��o(ͻ� ���7���ì\��2l���bX�℁�lF�]	
~ao.\C�k����|�i�^�Ax�6�װ���=Ȗ�������(Q��;��b�=�OcDb==�&|���BY��l��=5;}{2�/z�`6X��3
�v�v-}�	mpҭ���^���b��v݋N��������;B���Y���� ��@s'R�Dd�-$#�0��(Q��;��b�=��?njS���A���B���A�\>W�/Z��B���[@���[��QPw��r|��߇(���м	I���������)��H�'J!0��A�6x���9#�n9'��r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�^܊@3+'�tL�c>��*�^��o�������|I~�I����͵De��2Q�����ݟ���O�͛PA,q���R�*ؕ��A�\>W�/Z���N+~�{-M�O��~�X������<�N������ᴶ;R�������\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[���Г�D�i�^�Ax�`Vk���|�zYק�̒�H��@!�#-�[ҭ��;�fIx�x̛uBq����}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-��|��������2���t����)L��b��~���"~6���aq��yx6�n)_���fx'v�ao.\C�k�Ǆ}�tF�W�1'����
39 ;��x}��q���3B��*w��5 ���LIf��T1�"��z3�:��c��%2���ʏ!����>2{�}����q�rX�]��C`e�n
V~$c��X	��MUt��!v6�RMS��e�^�e�/��r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�^܊@3+'�tL��ɟ���c*^��o�������|I~�I����uY�0��f������C;�,]�eT٠�Y�����|O�\�+�q�� 6x�@�޵B�
�#L�tD:��@�JﾥI��P3�lWD�����`���9�#�PA��n�{��l[hbvk~�#x��d2)#^&|���BY��l��=5;�D�A�'�Go��<e�Y��%,��7n��dY$Ǯ]s������&{�zYa�w�X{��̱�4z�Tqn�}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-��|��������2���t�h�N#�Ǐ��b��~���"~6���aq��yx6�n)_���fx'v�ao.\C�k�Ǆ}�tF�W�1'����
3�м�1#���q���3B��*w��5 ���LI�0?2�U�w��r|��߇(���л���.Ȃb�����V�I�e!��nH�W�t<wN����#��%�T�s Wd2uUrG��Da��S�SI�Qq��D�|�J���t��B�F�4"��B�*�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��N���8@�we ��g庌NA(fۉ���$,��F܂d�ۤ�m�>!�����1���A�\>W�/Z��B���[@���[��QPw��r|��߇(���м	I���������)��H�'J!0��A�6x��箃R�@زB�R���>_PI��d���ˎ]":V�U=@:�-�X��WG ���b��1L��A�6x��>�TBΡ7W�FA��mӡ���<K�#�f�D��&{�zYa��K�SkS��9��IM� I0���ԏ4tv�l�ν�s��U;46��R��O+'�tL��tba��U�Ut�\�|��������2���tԷ���t���3D�� <@��fG�H�*x�߀�q��Nʉ�(Q��;��b�=���B����1��r�.Gb�TG|�w�<���\QqM��X�~ ӫ/��mbФ�حE�\�G����Y���� ��@s'R�gXk����$G����N�����,eS=�oA��$�J݃����t������~�j5r�n0��+c�wwH$��X����)ͶG�q�5Ւ��(�m��Xjۙ�)��s���d�7�X xO����B�}�t�ё�F�]	
~ao.\C�k�Eg����0�5ߧE4��J�1���Օ��/�����aq�z�1[FQ�񺗮���z��K	p�ၚI���ln�λ����#<x�5����`Ko����Ȑs(�"�H���o��qo�:���$��Xo�V�W'D�Fy�_�-9�#�ڊ<?@��[	J��;�P4ǲ �|7��K4�+Fb%��C�h,%I��t}�=Ll�����,۽��Z�A������sQ[��"5�o٥v�I�vv<Lq{�f��a��2�u|�&l�����B͗V�5"Y}��&YG�$���g]�
m�ٜgL��i8`DQ��Z�d���M0~�J�����`N�z��1��M��If�Nd+l�Yҽ֗�B�V^� ��u��.t���M�.ѯ�>!�&���Ԟ-zq�)����'�Q4�*�N���m�R����8�n��a����F��}/9�h�T�QN�~lAXg$���p6�ߏ�U�ڴ���e�ġ/���~���Ԟ-zqD7��@h�����HZ��Y��)�?Z����b`��Z�Ll����i��:
�����+�v>6륷	��h�����	�vI0���ԏ�.fOe	Ln��S�W�כJϾ�ig()��ikp���H����Q#�?���;���N���(���Y�P	dU�1�%WJo��_�n�To�[�C��-��JHn��z��c�Bo��\�H��/Sg�w��'o�7�C�j1�����	�v6������1�R+-h]GZEh5���'n�^0o��Ha뮩J��GZ>.�0��rF�,fX��"5�o٥�rv8E�m:��>��� ӫ/��m����^{�HUv�׿eJ�f�A�|��&p�!o躤/؞�{��X�i�R�ռ�����|II���XԮ�%Ah�%4
>��XP���v�c��Q��"��0��C��-���.x�1斄]��9�u�L��*����~���倽p�'ǒ�ƃ�b�7�*�7`����M�Z���	l0��F��j�
����uK�r�&U������G|M���9�����8�>r&���c
� ��Ces"��)Эb��v݋N�������8j�4�I��'���7=����2PW�uD} ���3�ҺIÙ=�H��M����A�m�(�J�>��?�4��icY�G�˱�ߓC娤l��&d�X0���b9���'$�HυL�r�&U������G|M���o:��
��/؞�{���yu�*����^��y6�T���1���
[/��̟vzL͊�q���z��e��Ɛg)x�D�����X���55+��>͌4s+�ny���.�R4��������p@�7�9�C��!�CA( ����_�s꘤�ID�4o�2d�F�����a�ɒ,��N��g()��ikp���H���j�(H(�<om��c�`�����Ћ�l�T��B{�LϬ9{vw��~JuAx��-r��|ڑ�H���o���� ��j�o]�����/� �UR0�}D�)x�?{���x.�KnqM�����ġ��,�Z�b8�i-EWA8���l��))�*���<�Hr�Ki0j@$��U� ���_����P%t+��m�yo�7�%p��.�%m�.�#7D��qs"�kV���"�V�p-�8m�1�}�0&�ܫ `A��~E�x-��)0l���D	��U�G�	�Q���e��OA B���]!�e�����c��%$Z'RpW��eB�1V�n�~%˼g��� ��"D�+�dI��'�V�0L��{�*���<�Hr�K���Z���؅��FJ����6��S3�ߟ{���剑bwZ_;��B{�LϬ9{vw��~���oaM)V���"�V
�Z?�3�����g��� ��"�F�*���_���D	��U�G�	�Q���e��OA B���]!�e�����c��%$Z'RpV�0L��{�7ȁ�$6C��[����7�4����5�%��/q||�S�
���N�@E�V)�jP|B�1i!�_a��zL͊�q���i�C�% L����6���$J*�Rs�08�b(���os0c��ZLN�	��2�V�a���%BJ�g
��4�d�cX~|�Ḏp�+�w��b9���JI�5r{�Ż�ay�Ȇ^���x�k]m��Zx�.���E� )�&p݉�,��}p�m~|����� �ܰ�a\Y����+���LQ��b9������U.6��̞��>��3
�v�v-}�	mp@�s�p���.ᬵy���"�n��T̞��>�h�5,Wlr�r%)cA>4h`�1�/o���͌4s+�ny��� �ܰ�a\Y���[C�W�v/��1h=��d����zL͊�q��C.W26K�~BvGޣkQ�A���ۖ��S�<Ԣ�E,�J�|R�ZLN�	��e�]#TjI��'�����7���{r��I`1R�Jʡ\��ԙ��'n�^0o��y�v�1�a-���7a
��r�^^��<E�{hY����r�?�o>�3�lrև�"�GI$��ǂcY�~�s<��MR�ɧ�	tc&�j��1�a-���7a
��r��L;Л��|#9����$�+�,�|��{�r1��j��Mشˇ&�,�>п�p=	�˳͠m�xW��9u$d9��}ϔ��J�s���
�k��!a�tc�&ck��};l�-���L;Л��|#9���hY����r�;*�}Ւ�~ܔp�l
d�o�R�N:��,��g�7�s<��MR�������c�A�L'��!�a��5�%]���a(􆿳��?ƾ�؀qjZ��H@H�֦g�㎏qló��|�����V��ߝD9�{��灊�O�i���Z鎬�������(���o���ia���lC��U�T�\ �͉��45�c���� �k{�� ��*ܑe�W����n�4�Z��g�p��;*�}Ւ�~ܔp�l
d
�3�x�.H����8�
{m�����`y���=�G�
>���B�5{kb���n;*�}Ւ�~ܔp�l
d�o�R�GI$��ǂcY�~�ː<���go^3��V��iO��]��A3�(N��㎏qlóm]�$I��I��'�ct�:��RE�QS����>�b9���S�nU�&u������u��U|<��⏇���;�z*���Be�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cULjaGkƊ~F˯�+)�F�������T�\ ��rD��+-�0�)7����|!p�f���CP����(��Qn���ɡAdk,I������/�|��(`��ү/�O'�=�1#��Z�����XP��ȇ3
�v�v-}�	mp@�s�p���.ᬵy��H0@&ɡ��r�&U���0��PWw%Ǧ6�ى��(`��ү/�O'�=���AJ����������[�x�X���+���LQ��b9������p@� ���t��f���j���M�I�h�
MQ9�F����RY��݁.�qO�.= ���V�6IWJE�r���秹�3I^�v�%j���x�;��ԁ[�x�X���+���LQ���"X��[�6�_��f�\7vm�܉��J���e͉�Xk��%�x<�<^r�m�����ч��M(���z�R<�����á�~O�2ZD")��7ǉ �Ş(�/�K^b���n�J���JT؛>�a�W+`�x�oP��@t�&�e�5
�������N�@E�V!:忴�n���o�4|Z�j��?�N�@E�V����P3��:`D�h�#�*"v%)��2�����_�f��ޢ1�a-���7a
��r�2ZD")��7ǉ �Ş(�/�K^b�����4��^��\i�@^7&ģM�'n�^0o�<:�W�_ĝ�gjo7�2}�<��b��*�ٓ���S���`�����ϼ	�
\#ȕ������T<�9�|Z�j��?�N�@E�V)�jP|B�1*)�)q	�cY�~�"���ʷ��m����-@��F~*7���&�_<���B�)���E�hxǉ �Ş(�/�K^b��6&��^�<%̚K"��+Bo�A;h�F#"�G����o���*ٝ�/�K^b�;��	+���f��b�������z��d>�Sg��%&I0���ԏ�.fOe	:`D�h�#�*"v%)��2������b��v݋N������&�K�+��&��Y=�ĵ�"xC���]/~�l#ng()��ik�:Q�l���˳͠m�xW��-#��k �&[k=[hbvk~�#x���D�#3�/��=6�s���"[��g�7���ìk���͖w7e�\��� �Ĩ�z=R\�U_�+XمL���BN�.ᬵy�໼�-xZ{S\7vm�܉��`~�ߪ ��e��R���x����ٓ�عk�|�,
������|�FIsŭf�ҿG�p�PR��{�&�8���/��Î+,�C��<�v�(|���;�ߎ=�$�Э%{�;���;�L���9�D_�3���U_�+X�M��w��k��T9s*��ԜF��Y��^��_*p��nk�r��VYW\y]/�qF+Yi=��o�IÙ=�Hw¹��<d���	fd��Q�b��3R�^Ƒ���P4ǲ p\匔'������^[_�e��IÙ=�H��M���o�G�m�?S>g�G�eI��'���z3�:��c��%-g?���ųJHn��z�F�x�aK�k�����9�%DC�2q�+��Ћ�l�T�����.��4�F1����������JHn��z�>�ack���A�;�֋`N(��/沄�J��CK8�Kj��#��'��wb�*ܑe�W����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85��p#�j\1�Z���=��L;Л�������� ^��y�C�ܨ�S��)�c�V�v�#ȫV�
nF�̒�Px<Eϛ�&�'�u��.t������� �\Yy���L�XuU���-��S�v�K�4R ��N��>�+���A[��E};l�-�����ɒ��JHn��z�;ӈD}tKD�Ɛg)x�D�����X�?bE��t�Y_�n�To�[�C��-���I����Ɖ�Uʚ7�ܩ�.fOe	3Y'zd��I))����A�m�( Ւ�XNQ�>-�W���M��2�B���l�2��Fm��b9�����e��_��I))����A�m�(�O&��܀6������1�R+-h]��!��q�F����j&|���BY��l��=5;N�����O�%��/q|��n�v��;^��ԭ�ʿ3��pApzL͊�q��#��}�y�,��Sq'�4bj���q}�`��@I��'�Π��yGb�-g?���ųJHn��z�F�x�aK�k��� ����H�ʱˡ5����o�إ����	`��nH�W��ө�\�5����`K�z~~�Y_"R�W�u+Yi=��o�IÙ=�H�R���}��M�+�e0��Tqmp�AJ�e�$�,W��+�Ds�`��=i���Կ,��_Vl�A.;��L�O����K���Jҡ:p����f������k��p����=bzx@�%Es �\Yy�����=:VFqB��R�ѵ�Th�f7��h��Ǝ>c�����eR�ʨ��_�\G��4�	B45��|49v!S�!-�+_d9��n��f�NDM�99���|1ugW��ZK>1wIic�a�Ma�v]ר)F����kI��'����0/�e��9�S���ތ�1��\�vŁW�����+���LQ�ͧ� �+�7���_�\G�k�y'��a�#%G����I��'��i�_:�ܯH�MPq6.JHn��z����s1�Z���=�U�I�x�؋�$xC��<i*����\P���	Oe��-��f�V�0��yf�1�k�����E@�χ� C�)�8D��N}�E�{פ>�>��5�Y�w����c��F�?�w-�s��|ڛuC,hG�p�P�+a�7��͌4s+�ny�X�D��H�MPq6.JHn��z�%�,��CU���it	�TU����z~����.`Ϊ�/-T)x�?{���x.�Knq�]���7'����eR��x#2���p�����h��x�]�V���KD:�}����=8ν(I��'��c8?-+eN1#��Z�����XP��Ȩ/�W�,��?ׄ/�L��{9�%��Z�vN���zL͊�q��io2�&H��ݫ�Q�����6�Q�%�+2�Ax���r!uA�T�g�v��ёo��%��/q|�c$n�&l'�x�Tu'�yK�w��b9���������]3X����a�x��M�ݭ�~r}*И��&���nH�W��X��:�&$*rv�����zY�l�Ʊ�_�eD�I�V�zcj[�����eR���oꘁ`�%A��C1#��Z�����XP����o�7����������Z�<ͯ�G��R'),��`�"z��q��p�AJ�e�$) u3��u"�������M���R��ӟ-�K䁊��l7c�{���=�k2B]p3��\0�N�}�Ȉ���@�ln�~�.�p�2�zm�:3��Տ�L� $�3"���N�T<1(�d�����eiRK܃��hbvk~�#x��%��#��#���F��-��j��Ů���z����i���	�Ȟ���i!�_a��zL͊�q��@!���X�6%V�J��5����`K��=!ߎ�΂l��=5;e�_�TQ|ò���
��_������,�XM�����0i���|W;/g()��ikp���H���lʭ�i/�Yx�y�Zgl�D�YG�9V���"�V닂F�Ӥ�(��Jx4���N�JHn��z���7帘��m���z�Б�Ty��q)YϦ�7C�\�H��/Sg�w��'o����v�]�Uʚ7�ܩ�.fOe	��|�T������~RK܃��hbvk~�#xeayA���r�&U������G|M������1x �Mt��5�ء�Ch�1Ǥ �)�?�0��Y��W���U�dP_\G�7^2$S�6���f�_)fxg��pH���0�Ҋ@)�t�d�f�rЄzɳ�B��,��C-2�^���ij�IROgn�t���c�&�<�o��H�,>��*�:��I�}L������@���t����N@<����fRD�}a�/^�yQA��D,��f�x��r7�1�v�������bpQl��u�!�`�(i3"�,�>E���]�!����-ዧ�[d�x� �q��ُ<��%!�`�(i3"�,�>E���]�!��	Ǹ�y85��_�j^�I4��欱���j���w�:Ës�yb!��u፤.��.f�g�FQ���|*uN�wHZr��AR1<]Q�I����踫g(�r����*j�B3�&�#�vi3�|)sՀ�23
���v��Ŧc�ƇBHx\�'���Xw s4S�'�i��`�z���n�j�Q�c�_�����ʙ@E>*���ls�u°������R�wX��}�
�?�a���k�_g��������/y��g�'b�t	�U���C��O]r�<Uee�N�����z%$��h
P�%.^F�	��lC��U�T�\ ��i3�|)sՀ�23
����X%�(�ƇBHx\�'���Xw s4S�'�i��`�z��Y��)�?Z�����1�����NR�^Ƒ����"X��[�z�C���vے�(�i�p�� �&f��vA<UV$�����wY�{'%s�[�&B�踫g(�r�N�ǁ�f�TЏekZ�>5i�[r��5�%]���a(􆿳�f����DB}�
�?��:�,��mj�(�������Ր�z*���Be�2l��4��a��se�ξ���e�J�Pn\�pD��ZOUi3�|)sՀ2��2,��g�ܧ*y+k&v�IzZ鎬����
C��8q��f�kN�ı��U��+�Xa�H(�˕�&Ã�M�Ĉ��r�]@P�B��X��8���/�I����"�Oi9L�:,�۞��	����YLZ鎬����
C��8q��f�kN�ı��U��+�Xa�H(�˕o�`�_f>&�&i�"j���b7|#9���b!��u��N�!�`�(i3�􇃬Tk�H@H�֦g�㎏qló��@d��ץr�&U������G|M���t�2���B�D�F �(����Cb�\�V��7s�9���o��S8�(´W�w#�m��P���ݪ��°������R�wX����K�Q]���!E�r &
�$J�n`5�fK��0z�cUL�n����4����it	�TU����z~���ӯIJ ��`y���h}Nw���eZ���08:�}v����]�!��	Ǹ�y85��L�@��f����k��$a(􆿳���2����.\�#$�ÙA;��W���n`5�fK�\w��0]b!��u��չ���1�JS���$�q���U�h}Nw����;��[TM����z�Ji�y��Fp����f���,(���B���̴_��EI?�R��n��am�Za(􆿳���Qs���Ѕ�HN9��c�fi�d� ��^�:AԢ�a\��F�dH�Dj���G�Օ��qvdЧ^{�j����#oM������ݓ��E�S���%����g���hZxZ��j�
�iB{�Z�_�vW4��`��Q��ǺΕR��ӟ-�F`���G���`y����@����gGf���ѩj���m�7_Ņғ�vq�\[$Q��
�`�ю龤9>(�vgH����8�Ј�&��g3�g��U-�e5��e6²nx��hѧ�����n�۴1��r�.h�k��T9s*��ԜF����<	�'�K{xN��i>R��n�J>|�
#�`�^{��u�oD�|.�Tӏ�;��[TM���!����'�U��=+��K)zum��3A�)Oqy�&�CA�R�.��On~���=���q5�n!_���'F�7��"=���;�m�PV|7��'�b���b�Bϱ���w�K�̄�Bq���ZLN�	�����#oM�������׎o�|䖬n���!�`�(i3�d�o/�d��7���ìk���͖w7a&r"� L,pzl��a�T�n��a�I�T`��$��qgo�2}�<��b��Z1�i�a��ġ��,(��T�eȘ�Kⷠ/s�1��p� X���/�K^b�Mc��_����H?`��K�Qc]p�5�	�7�|�ةGy�ˆn����Sb".�f\�H��/Sg7��yY���k��VPI��DP֞ M��V!�D�n`5�fK��0z�cULjaGkƊ~F˯�+)�"j���b7|#9���b!��u�+�uB;y�������Y�{'%s���'����C�`�/�t�KV*�3?�|��T�5�d�,WT	W $V��8���/����,DY�O�~H@1"�,�>E���]�!���e��Ƥ����n9이J��sr�lғ�vq��/��j�3�T�\ ��i3�|)sՀ�)׺����e���b��d�٣���N N�S�qg2�K?\�2�q��n`5�fK�\w��0]b!��u�#� �,W�_�S�
ut�q���U��@����gG�0����Oid�w4ZxZ鎬������_�,��|[p2e�F;p�	�j}"K���rs�i����ej1W��Mw���1�Z���=�"j���b7�������˞�BxCeFJ5x�_S⏸[��!�`�(i3��lJ��튝�b�Bϱ��ᵉ3������d/h�5�G�G���M���X"�,�>E��P"G�wk�١��	;qBvGޣkQ�A���ۖ�k�V\���"X��[�����O/h�5�G�G
��7t��i"�,�>E��P"G�wk����Jg�|#9���!b/����Я��7�Ixi��z<}��\=%��I��'� ��k\�D�1d�Fv�x z�Jm]A�/�����`z��V�%��/q|Kǹ|���:��kdO������������]'ݪb:�B�eʣ͜��խ�~x�;i�?�rn^v��Y���0�ȷS�J���]6���b9���A��LE�Q���'��{ �=�%�,zG�m�yfÁ��/�ϟ�󓅅g()��ikp���H�����bK,��G?�R��nI4�p� ^�b��v݋N������<�bu�C�b�P�b� �I))����A�m�( G��+�a/�K��]Xgs	���C��	Բ�`J>����:ҹ���7�&k��F\�1�|��g}$�%�� �jPxT�l�ޠEnݡI|4�8�"�6�#vkɴ��F�=��� *�v��6
R:SwL���"�R��@L�_+H�]��Q١Ӿ�$/s�1��p�E����FAԢ�a\��F�dH��e@�N�] �v"��x�l�<Ң�8���/��Y�r�7"�*��9W�����zՠ�F��6��U,�(�)8���0y�	�C�u)�6�Օ��qvdЧ^{�jt��zh+�,�l��=5;.���������#oM|#9���7��"=���!��V�B���.V��:��^��[�@g�#�ڊ<?@�֫��XA��:K�e�>c�.A���]ߺ�`@��8�v�@����n9��wqMYxw���UӐl�L��M�,���	N^�U�}�g7�}�ξ���I��RhF���9���x�����,DU�m#j[ql�d_b�B�E`^n�&�
_�n�@/%{�;���$��dg0J�I4��欱���j�����0À�C���DP֞ �g��n%��gn�=4;J�F���A3�(N��㎏qló]�b)�L�uf�Nd+l�Yҽ֗�3���W
�����n9�����[m��3R�e��2����@�*ܑe�W����n�4�`t��D����M����A�m�(��ڽQ����M�q�Z���U&�Pֻ�I���I�����O�L��pa���c�SD釛-���>Tf�Nd+l�Yҽ֗�°������R�wX����K�Q�3R�e��Ӵ�"�6j��;٬sf.��$T�=�|��{�r�]#I�P�*�7`����M�Z���	��"X��[�z�C������N���c�v�_����J�����IhEUE�?�o>�R��}���N�ǁ�f�T��p_U
#�g��U-�e5��e6²]�N��&���3�L���'s{	�h�v1a{J�ޥp�rO�`�|��K�z�Q���l�N�����:��6}���8���/�a'�<� \�e�bn�m�±��m|�ժ�E�$��*�]u�W6��bS`�|��K�z2u?r���Y�G�˱�ߓC娤l���Mq&�������DzL�a����g{A�dha#4��������y� ��[�$��X�՚��l��H�/�n>�.-,��Sq'��_�H����K�Qɲ�cz���ł)w���m�±��m|�0ί�.���n`5�fK��0z�cUL�JJ�4(oW/S��8(�E���Kt�m���i�s���1�R�n� �}DG�M���f ���`y���pzl��a껎��YxP�B�>��֑xGV�2��."�z�����R���q�41&q^�`
�c��><�$N�w����H��4�d�cX~|�D̽��K=$r�8���/�a'�<� \��|�fL
��"'��l����C1zh�O�P\*=3� X���/�K^b��6&��^�<a'�<� \��|�fL
��"'��l������O���FW��n`5�fK��0z�cUL�JJ�4(oW/S��8(�E���Kt�m���i�s���1�R�n� �}DG�M���f ���`y���pzl��a껎��YxP���2�ę�u'b�'=�(�hU�AG��q��T��J�s���
�k��!a�tc�&ck��Wڭ��h�Ɛo�c�?EcD�=1]������R�wX����K�Qɲ�cz���Ӵ�"�6j��;٬sf.��$y�=N��"xC��-�T(u	M^ڐ��S���pzl��a�	�_��:��u���'b�'=�(J�}�֖�c���[�s�N�@E�V����P3���2��:�k�t��S�D�����X���*"��Z�w�l#���i���N���c�v�_����J����{0	�b<h�d�o/�d��7���ì�"����x,����a�/�n>�.-,��Sq'��_�H����K�Q�3R�e��Ӵ�"�6j��;٬sf.�r� F�3N$��qgo�2}�<��bl���>s�q?H^��2\'P�����M@�qX�Uu�T�˷Mq&�������DzL㡉�&�@�}�-��w��k]m���#�;�\���J���e͉�Xk�
̄?�90�ΩyO^~~���=���q5�nC�)�B�Hpzl��a�N��	�Ȓ�@{2귑���Ӗts�T�]�!��M8���	D%��_�ͅ��r�&U������G|M������{q����'6���;8=�g��U-�e,%�0g�����L���N�b�'BeoP�z�y��R<����z���踫g(�r�x�y�Zgl,�B۸�Qz��!"�����;�B{9��#.��"��J������-VL������ l�\�n!9�*q������_&���I�*���Wk0F-X	�4�u��u�s[T��n��؍ݓ��E�/������-Ӥ�v3Lp�6%Y�z��d>����C���ﵒ�v�{lGD�V�B	3i�\��׹��t�'jG+�$�H)}���/��C�x!�H�Ȟm�2GS���J���e͉�Xk[�[�O5��M�q�Z��1N����F������m"���g���Y�{'%s��.|Z���I7��-5��6��	���`y���pzl��a�)�O�=�}ҵaM�B��5��k���{|�rs�i�jf� l�Ǜ������CyW�f�tR�wX����K�Q�L�t��n',Mn�Va��W6��bS��A3�(N��㎏qló2u?r���Y�G�˱�ߓC娤l���Mq&���[�=�5x��j|�>�O��R���k�:A�	S�r��AR1<]Q�I����y�搲)���$:N�8.����6a'�<� \��y��`_��F�:F�,����};*�}Ւ�~ܔp�l
d�R�.��On~���=���q5�nC�)�B�H�
�CӞD�2��@N����B�m�=][e���w�<[a!�����QB�cG���*ܑe�W����n�4�{lGD�V�B	3i�\��׹��t�F��%{j��K�Q��������+:c���d�٣��c�A�L'��檆�R�wX����K�Q������0�� ��v�d�٣��c�A�L'��檆�R�wX����K�Q��6U(�<"�%�մ�d�٣��c�A�L'u�6949%t��R̕q���s���8���/�a'�<� \5�q{?za���{2��D�n`5�fK��0z�cUL�~�@�[���}�pIɽ�Jz_ꛨg��U-�e�_|�<���T�e�V����Q��uзq8�Ј'���Xwa'�<� \P���Ʃ85�k80��߯�k���{|ό���.���K�Q|��L�����Q]� _�rs�i�CЎ�����Ɛg)x�D�����X���iB��.8������5�e`��9��\VO��1��0����Gs�	d��0z�cUL�~�@�[���}�pIɽ�Jz_ꛨg��U-�e5��e6²���`���l� mr�m�ZsD��wό���.���K�Q$��Ly����:���@Sz��맆�q���U�pzl��a�o���
^���|6?����M����R'���Xw�j�7��	w��������΁In|��B�S��������B�D�F 6�W�.s��錛�%`��Q]� _�rs�i�ק)"�僁��{9�%��`0P� U.R�wX����K�Q�N�]�B���vE��nK݅�Y�{'%s��jb��:0X����A.�%A��C(Q6D����z�C���0��jOT�Ǹ���)/�~�T���]�n`5�fK�Q2�+�Yɳ
�CӞD��g:%���5�>�k��q�9k��q���U�;Ӭ8���o7@w�MS�sCLq�M�7��jqo�_h.\��<Z:uoZ��2����E�̜��W��)�mS)/�_����f�c\?kv�} o7@w�MSʋXr�$��2����E�̜��W�����5�锹,hy�̥͌!����$K�A��2�����z��I/r����=q����p��u���A)VUegrE�:���@ŋ��5�$�)=��r F�)tH�#�rU҃��~��b��T�Q5�T���@W�s���CL���-4�B��.��~r��9�c%y��dR-��SBB$�W%�S�ts�'����o���u�X�m��{��N:��")ݝOv%6�!	��1��yt(���+c�(Yw�A��v������m�Z���ё5<w�⽒���M����A�m�(��D׉��h��$1&O�Md�sω��F���1���T�}ɻY~�y�����[�T���Ӫ!��˼�v��j��gn�=4�D-'��7�q����5^����rh��,��G���۵z ��gn�=4�D-'��7�q����
�DB�%�$����Od-@��F~*7���&�_$� %7�zf	�$NT�I���I�����O!ݨ���0���º�>:��_
�u��Yx�I���I�����OeU���(�CK{D�sss2����`�|��K�z>���@]Ps_*�GqW�w��fD�l����lѣ͂WL�!�]�5����V��F���1���T�}ɻY~�y�����[�]9�(b����˼�v��j��gn�=4�D-'��7�q����5^����r���o���F��!���Dڋ��mhcA��짦���O�ʦ
���c�v�_����J����肥�J�p�0u�xs�&q^�`
�c��><�$("�P��_��3�.�J�s�xV��8���&�@�}7�q��J��v1a{J�?��кDO�YN
��)e�n�ߢ���8p���uAԢ�a\�DW��E��q��u���'b�'=�(J�}�֖����%:��.����7���{r��f���꜅�R��ӟ-��>#qBK"6j�"Hs!�pL_�g��L�*��6��@��XL��a��������+��T����oGo�Z�������/�)��ɖ`ۺ������Xc�F�������ϲ�>e��>��0��E|�,VK�5��&q^�`
�c��><�$���E������Kp&�w�%b��G�w�Iſ�Κes��O�h�S{�5��lW0�c4�j
Թ��~��q����U���*'<���h�wIk�� `A��~E[q����*��b�&z|X�L-�.nN7� m[��G�Hl�W�uXSr���K�H~S{xv�D-!�͉���ڃ�"��
!�7��}���3r�dv��oTN֢&@��&̲�2�!��0��"��S8�TkF�����3�L���'s{	�h�v1a{J�z@�q�H�[�t��#���n�|����Y�{'%s���F���gn�=4�4�	���WdM4@���X/H=��q��G8��5aU0Q0�wqMYxw�R����Όꢤ�Ogf$n�L��4�g��n%��gn�=4�~�����9+����qM�o��8+�)�y���mcl�y0q���Q�L���\�LtF�/�X�h�9�2Rr&��Ih�	�;�6�l!x���M���R��ӟ-�F���ˏ��Z��zf	�$NT�I���I���C1zh���\v2:R������S�_
�u��Yx�I���I���C1zh�6���Q,|y�����Y���ǡ�C�a\Y����+���LQ�s�xV��8���&�@�}7�q��J��v1a{J��ש�
�~��,\���ӟ�X���&�@�}7�q��J��v1a{J��>�_��� �U�N;k��!a�tc�&ck���>#qBK"6j�"Hs���ٚj�ώ ���]q޼��B�p,�f�s�G�6�l!x���M���R��ӟ-���4�&����Z��zf	�$NT�I���I���C1zh���\v2:R8�dEm7�w�kkr�I�;(�\��8p���uAԢ�a\�DW��E��q�����C��֑xGV�eU���(�͊����ss2����`�|��K�z˦9��iժG�p�P���ً ��3R�e��Ӵ�"�6j��;٬sf.��ǞZ߻����zk2�����n�۴�.�<Mm1���P�|T����E�E��3�L����e�eV�M�z$��P�^�6�V���l�p�H1�a-���7a
��r�$Dc~4�A)�V��/�c����sL]~цt�U(i�z��Ά�A�C�	~�)��u�X�t����r9m��+���J q�v����6��w�1Lſ�ZO&����S���� "5�]h�' L� U��֜��3�=���Q{�1�a-���7a
��r�b��j��<�I7��-5l*���T�I7��-5��5Z�����L��c⳯���Eu��oŹQI�~�џ0I� X�1� �����b@c{{��
J�~���.����7�*���<�Hr�`�_��QA3e��q���)��j)yc�n�.�_�t�H2v���Q�[��C���������a����"�$k��,�:�N�*�x���D)��g�%Y��̗0z�cULj� 1ɡ��&�@�}�-��w��k]m��>=!=�"���Mڷ�l��)��'���Xw�j�7���3R�e��Ӵ�"�6j��;٬sf.�B'=�:�,�y&�/S!��4_���QR�Xe����;���/�kI��Aġ��������[m��3R�e���V!8P�24%6� �7��)Q�XI��J�)��yf���x�M�g�������*[UxG��
�	?�<�a�/!O���������T5��t�\��ot[�W��Vg��{�����$�(��n� ׵����:�#T�a��p��x+6���Z��~����p7A�SW���)�aO�j��&����KS'�*p��0���!�|~�X��˓"��0��HXC/���eV�
��e,OL���t�b�hO�^+���\5؃a~y=�,����ێ_ϞB �'@v
@�1�Xׅ�LN��A|���]}����xT���b�c�r�{jFKL���:�G�h�� oj�VO����+���������᥼�5�/͆�꺖Z(��:�l�5�����xn�|������Y��#�¡�kU�%Rd�B���^��5��f�
�7�gŢ���ᣊ��f�T��nxq�� +@���))P�����X�C�HC�|��dq9%��9.7g�t���<���/�3��Ay&<y�;��|B����N���h_�zG6�o8:4�I���c�90��c��qq�KX��ik���`+iYb"Όd)��i?|	.�4��s��Z���.TE�g�������(ӈ��� �3�c`��0��₎���Ȝx�5W ��̫(>��o��X[�QB���X��WG ��i?|	.�4��s��Z���.Tv{��lw	����,Ǣ�Пe���;u�4�J��x(�i��/Rh�x#�L_�(D{ͬ�y��IX0F�M�^����'�֫��XA|>���)��뮗�w�ތ4�7�K�Š=ԕD��6c��wV��߬�F�<�t�W(@M�(fw���'�̗������k2m�;��|BG�a�����C1zh{A�dha#4��������o�^Һ�^E4+у��b�Bϱ��3R�e��ł)w���m�±��m|J�}�֖���J�_��e����7���{r���i���A�* ^��\�v'b�'=�(�ժ�E�$��*�]u*+l^�V
h��,��G���۵z ��gn�=4�4�	���WdM4@��&����˶�6�>��ʬ���7���{r���i���A�@[�_zβr��o��SO�W,�P &�\iT�������܏g��L�*����`w
��Օ��qvdЧ^{�jM|�"D^���\�}6��~p�=�J����6x�F�-LU����{����J�^��4br�����w�����P�<�F}���V6��Q��&i��N�N-��;��M�z$��P�^�6�V���l�p�H1�a-���7a
��r�$Dc~4�A)�V��/�����;٬sf.�#@�Q¢�r}l��L�e�+S��2v�C�|J3J��$5w����k��뗁��cA��짦���O�ʦ
���c�v�J��sr�l�k]m��+qO1U��#_"`��Rss2����`�|��K�z˦9��iժG�p�P��c� V��	��yv�ʯʗ�bu�r��c7�
W���ݤ�E��p��4#h���C�m�t�T�.�p�ݷ���1Kޑ�l��'�.ᬵy��̒�R�K!����� hbvk~�#xXX�dPh(??�d���&���xBS1Or}l��L�_�Źz=+��T����oGo�Z�������/�)��ɖ`ۺ����L3�v-Z�^Q;�im����n��+ԑF�r�f�t_��/���-@��F~*7���&�_�}�����*�	s��NU��֜��3�F�7��Y�
�cc�V��ģ��N�/�B{�o
�@�Ce�<�`:�(	�����Q��K�g� ,�,jsUD������]��#�w�uIf�d�Oi��5K^�}M,�d��T��ޔhNVBN��
�5K�ƠX�L-�.n��B*T��� �8� t����$�¿DĢ�WZ��b������t��˳S�=L���Y'B�ɏ��]�!��	Ǹ�y85��*�Զ�m�±��m|�ժ�E�$��*�]uz�|W[?����~�ܾ~�X����Z鎬�������(����n17 �̿WdM4@�6x�F�-LU����{����8B���=�17�
�5aU0Q0�wqMYxw�)eUȯ���3J�~{������U��U�%
�bJ�ڣ.�����2�������E�i�5t�&��f}�~�cj�:1G0���oC�����8y����>�'~�1`u_=3O��H��b��+�+:�<�]�Ե�/��}&l�V��	��y���"��l5uS��~ �4���ګ.�0$��*�]u��l��'�.ᬵy��h��9h$�p���I�G|L��v�8:�y��D;��|BASf�<M��=�^�36�o8:4�I���c�90��j��e��0h�5e�ʙ�fZj:� ?V�)��a-6�Da�L�t��n#�%��>�h0Z�W�dN�<@Iv��nt=:ྵp�!����0��₎���Ȝx�5W ��̫(��a-6�Da���L�nM?��y�Q�(�r4���g��n%�)eUȯ�����J�^�R�Xe�������(2��y���<�K�p�-a�D͢q��`�L�5ߧE4�������`05�N���ȵ���m1�H���W�w��fD�'��m�A��d����x�C�����^���O �I�<^&!!HY$2:rvB3�c�}�C?����2N!�y{+_��F�:F����>�]/��=�~�1�W���h*
��#����[mߍ�C*��y���<�K��D12��G"��y"�6��ޅ7�=w�I��RhF��j���W���?�d���&�^�n��Uh��i��z����>�v{��lw	����,ǢL�E��<U&���8V��	��y�����'�s�I���Io��]%�TƮ�����[f�Nd+l�Yҽ֗�,�3�YG�^���\�}R�Xe�������(2���M���)�O�=�}ҵaM�B��5���p];\�;��|B%����$x��ڥS�V��	��yʄ��]C���X�C�HC�|��dq9%��9.7g����'.�ڨV����>�q&.&οib��0�>%��l��`�9:tq܃�KK&P�3�gTn����v�٦_��s�֙�;o7�<��j|�>�Op�Ńۗ}:)�O�=�}���N|�H�e�8�m
�X��5�fFG�j|�>�O򏇱�{�� ,��rQJ�ڣ.�����7x%p�|�+��?�d���&�J� 䋶�a���hJ�����R�/c��/{j��+�7�����?�d���&�D�w#p\5��m�Z�S?Ϳ�IK��`���-�
�s$�����Kӡ�S����		*O�J��i-h�(���b��b���*.埲�<������׉�	.�fS��X0\�^y�S&���=H~3�A�Â�v���ua�n�|ò���
��_�����pJ��y��/��^��:I0���ԏ�.fOe	U�f���n]�zP�w:Ec�[�p(	��e
��+�)�4B-���4R�Xe����ɲ�cz���v{��lw	�c�}�C�ǹւsr⍍N� ��"��������L}O��Q��nY�^䰃���,h��z�[��D��bt��N&ڸ��Fp����
Ո�C�hk��Y��A�m�(�RB���
��\�� ӫ/��m2���K��֌I�<�������|I�ݱHه��;��|B�cx����wZ��,x��C��7��<hjY탌������-���=a���iy8�b]�l���� ���B��[Y�QV�LC�5��}a��n�
�a8Xs�'�����q��9gc��@�Y���b�D4�\:����ϥ��W�Nʆ'��b���4�D�X��7��=Ŗ���8{��鄷�)p<3_�έXt#+sq����1�<��3��iie��!����m�3�% ޕ��Y �Y���m�jV{�������P�R�ӚO2@������Jtŉ��n���trq<�v!����W�ID5nQ�rV�sT�4�;��|B�7e����_��z3�:��c��%)���;��q3��+���-��Rއ�j|�>�O5X�nd������'�u� ����a���wqMYxwt�"߉�f&#p� ���N^�Yإ"i��V��	��y�+���jt�J�h�Iz���W��-��8PWa�X�w�.ᬵy��z�g>�HW�w��fD��dRPZ<�f������C;�,]�eT�?�d���&�Tc44�.������m"J�$��F΋�g��n%��gn�=4��Н�H	���0Exp��=���+.���!}�~�3��-�i�^�Ax�뀊��TU�?�d���&�@�n7�d��}��R�Xe����d�鳪:��X�m��{� �;Y��5b���t��P��M��%LS�����q�z8�2����v#�J�G˥��	�ώ ���]q&^�T ����Օ��qvdЧ^{�jmWᅫw�^���\�}ɲ�cz���Ӵ�"�6j��;٬sf.�����S`�^E4+у��b�Bϱ�ɲ�cz���Ӵ�"�6j��;٬sf.��w�b���k��!a�tc�&ck��Wڭ��h�Ɛo�c�?EcD�=1]M����_���|��
�|u='�c�-��;��F��zF�ۗ��ʼ��R(F}���V6��a[a��|u='�c�-��;����W�O�힬���7���{r���x�] %� /s��EB�w���%���ց���=E�S�Ӽ�26j�"Hs���ٚj�ώ ���]q�bfb��@_�bu�r&^�T ����Օ��qvdЧ^{�jM|�"D^���\�}ɲ�cz���Ӵ�"�6j��;٬sf.�����S`���zk2��������;���]�F}���V6��a[a��|u='�c�a����g��Z]��-@��F~*7���&�_5�NS�x�r�r%)cAk�Ղ����Y-��V��k�	�"�kϕ=��8�%<}���"'��l����C1zh_��N�\Y
�P�DQ��w�kkr�I.�rm��6�,\���ӟ�XC��(3���-��w��k]m����ǡ�C�a\Y���[C�W�v/��1h=��]�V/}�j��4�d�cX~|�D́.�.����|�+��?�d���&��$ͯ��A_���qmǵ�zb����2�ę�u'b�'=�(@�|6��]̷_��yC��S8�TkF����#�(�>^�l��e�eV�F��zF�ۗ�Q��L�
ɴ��z�D-'��7�q����������]�!��	Ǹ�y85��m�AD���"'��l����C1zh_��N�\Y�����pܬ������@�[��(����5���ռ�j����)w�n��ukh�)�_��,\ަ�It��+g[�b�ӝ5�T�w�%b��Gv����Y���a\Y����+���LQ���ll��4�(�hF�w���a\Y������bPv������Kp&�w�%b��G�w�Iſ�Κes��O�h�S{�5��lW0�c4�j
Թ��~��q����U���*'<���h�wIk�� `A��~E[q����*��b�&z|X�L-�.nN7� m[��G�Hl�W�uXSr���K�H~S{xv�D-!�͉���ڃ�"��
!�7��}���3r�dv��oTN�A>�''B�ɏ绎��YxP�B�>��֑xGV��Y�ٺ�rc�x�	��)'΍���>��[�s���J��sr�l�k]m��`m,�y���[b�0<��U�%
�bȷ��>m��=PRpY.[����{�j%a}�C}��VӁa���`�=���Aɀ��R|�`�s�lo���I��
�[��b=��|�)՜�4�vIn�����L�r/.�ij8��T|ڭ�F�\g�G!@)c�"j�D�)�c�}�C����R�Xe����NL��i�i��5Υ�ZahcZ�lF��p�Nģ�Z�4��6�zy�Vނ�L>.Gz�k$VQ}�!9�!4.'@�q��������0�e�҄��_U�C�s�6s�uƆ�!Q0�U��q�����O����2!�Aͧ�z��|m�Ř�/5���V�� /g�!���2(�4�D�5��rL���oy�{���;J+���Q4� 
A��X(�%{�����a��;�-mO���RLT���W��'0���5�� �Ֆi�8�oQk8�i�ѝ`D�c���*�9��0,;��[���j)�qzB&�|�dN��"��z��|m�?9&;���h��v��:m��F[ �4�Rkj}kqF��ہG1��^���fU�ZQϱ$Z�n���/�GW������)��n�V�����aǺ�#6M0�
F���^�����\;��~��M���s�A�j��@A�0n��cL�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��"Jc�l�!H��R��M��gq� �ɰ����Mp��Q�V��&��C5YD�H*�r�wl�({�x���	R�N~)�jm�w���i���Z��FkH�������h	�(����5���&<˴m�TJ	V�+�PM�^-q�x�l��1:�N�*�x���N�4���f�����Q�_f�Nd+l�Yҽ֗��k�+9=�]V�H7'�R�^Ƒ���)ύ^��R�^Ƒ��f�?ǉ�=�m�n���֣��n��ݜt���,\ͨ܉p����O,8�ݚ�Н�bs��2[������	�;�ݚ�Н�0q���Q�L��
�:qEp3?���*�YmC,igu?V��j�c<�s����	��7��u���/	�C\�2x���?V��j�c�?�#B,��	��7���=��ծœ��K����f�?ǉ�=2W���R0C7z���.��.f���T��M5��s������>��>hߵ�V��rU�w�⽒���M����A�m�(��D׉��h�#g�k��r��18�� TF��&~����ww¹��<d���lC��U�T�\ ��;��|B����=���p�� �&SfzF�.���tAC�����[m��3R�e��,z*ը����u���"6J���_��ocm����$Ȣ	!��.���� _>��>0i��.��J�������^�d�����w�>f��8�Dw]r���|�|P8}Ά�ud�H�A�m�(*��l�- ��pg^���W^G�2y���H�V���b�?C�F�.��.f�Cz瀿3�z���]�D�)�O�=�}���N|�H�ejxL��Ƅْ�k&N���g:%���5�>�k�_���(&�c����7Q{��̯Ǹ���)/04K��%�&n�i��V��yRf.ܸ���=���G����*�7`����M�Z���	(@��,1����Ѹ�Z{}t�\mc�#g�k��7�_�ܦ��X%�(�!g�lu/����t��P��M��%LS��b���jp��0�| ��p�-a�D͢?�d���&��bya�C��<^&!!HY��w���V��	��y�� �P�qN�h���w3&�4w�d��˩���.p!�'���4��Ǳ߁Ĉ��r�]@Oz)G�F�C�T�\ ��;��|B����=��F��׿]�v����D�ه4�tZz_nÑ2hꬺ��1��NjX�U�6j�"Hs?�Jy��{Q/�C�#>��G�Ȧj�E��g�Hb�t]�<Lz�����=�<��̀��unЅ����D5�|أͽgF"?f�Nd+l�Yҽ֗�,�3�YG�^���\�}GP��_&?Wcv�mAvWދ�qc:ct�:��RE��W��_��MM
��,=?�d���&�����x������v
6ڑ�I����<�W?�I��RhF��U>V%`�~��POۭ�٤.��.f�Cz瀿3�V���!�F?��G�Ȧj�rZ�0m�\�n�8�Z�Ѽ�;%4fC�6j�"Hs�2�p��΂�j�|JK
��ݚ�Н�Z��E��3?�d���&�o3F�ȧe��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI��ߎ�x}�IUr��Ӱ8��oZ<8�w\�PPOi�<ՐW��K1Y-r�EHd
0Ki�|2;$�J��7�OT�,��7=����2PW�uD}qb	��G��	i5Ɨ�}�IUr���v ���\{a���k�_K�ǟ
��)@[�_zβrꢯ�wv��QX�mR�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�wP-�H1�m��d�7��dt�{��!�r��I6�qf���?v�q�2�_:��p\I��� �W�G��!?�d���&�db�\EXP-7�vqq��I�?g�f��r�F�5��I^ξ��ݴg��S�ZC#fr�L��ϸ��#|S������3[�u8��p�ϵ�DE�U����L��g�e�J�Pn\�6^M����!�`�(i3������ET�zn�x'��݁.�q�0��E|�,�k�+9=�r'Z1p8 1���H-�`��E�ݦ\�t!�ǿyXAm�,���9^-���2��̪U��֜��3�kޮ��R�^Ƒ��WP�^:J�_���9�x&_FA"���)O�r�h5KQOڜ2��,�9�i9^��
��WZj:�Mpp�}�(�-l̜	H��d˹�40<~I�~�џ0I� X�1��kޮ��g��� ��"aJ �!,|�8��5ǛHO��E��������~G����EX��dC$,\ͨ܉p����O,8�ݚ�Н�K�\7}�W,:S�.?<N��	�Ȓ�@{2귑�7��m�K�!�`�(i3+�uB;y�e����'�N��(���K�!�`�(i3I��
�[��b=��y��j��k����U{8�C,0�?��ʉ��%>�rG�<�]�Ե��M0?n����)7����F�p�䘶'�,0��.b|��Aam�oT%Und�/n�-�6��Oa���G�usas��1�P&R�|S���?d�bYގEV��2܌��o#��V'U4��\w��˪?�-e�J�Pn\�pD��ZOU_��s�֙R���Bk�d9�Z�y�6H�S���BvWދ�qc:��S� ?�0��E|�,H��q�/���˚����Z�ם�.J7h��C�x!�H��Ex4*+�� m��DKY���k]m�����|f��I�{�P�՜���,�ǰ��������2܌���!��g�9��,Y�����9C��K�J���֏^�M;�¬pX��D�P�E6�k��q��־�W+��W�V;Ƙd�d��]���DKY��,�۞��	�>�A0_�|}�	76�&�;��|B!�{I�l��ԵW��;_��8W�w��fDbYގEV��2܌�xуr�w�R���y�A[�;��%���*�'IZƀ$�ֶ{�ӱ���9��;�R���5���T�}�@��'	�?��[�-���^�ߗ/�h.��t����~,�046dr����,�ǰ�X�t�q���Ù�?��	`��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��N�b�bq���Z�N�;�{W�5�St�IM˶I�?g�f�ja1�n�[�ެT�Z¤��I^��?�;��XC&��z lc�x�l��1:�N�*�x^�R@Κ�2���ei�&8�,�뼥<7.���nH�W�f�?ǉ�=K�|q��=H��6���,���eFz�p���,���<ͯ�G��R'),��`�ce|O�|�:(�I~�����h�Q7!�`�(i3����8��]V�H7'�R�^Ƒ��!�`�(i3�F�7��Y~s���6�����{,[�=·j�U��֜��3�&8�,�ݕ����׋�es��O'���OY3׿j�h�<�������i�״��/^l1�Z���=�,���9^-�VkLs��dJR�^Ƒ���X;p`����0/�e��9�SW�Ty��5������[��C��!�`�(i3�
!�7��}���3r��+qѭ�+g[���|��p�S�o@�����	�;��=����t�7��r�=H��bf�?ǉ�=�չ�Ad���c�����:��IK��<?KYC'v�����6Y����$�g�ܧ*y�?�+�p!ЈH����@�/�MC7z���N���q�0){\���Z!>���j�3���0��ĥ7��A@�r$p!!v*!��o���sp%'�|]0��؎l��%-���'��D��$L���G�+��%�k<�6��w�
=�2����޴�ik]�O��Z�l�X� �Ĭ1�e����:�ԑ�*V�D2U4��\w��˪?�-C
2��>�q;Rm�5�O�%E#P1h#��x�3>�G5��,vQQA�q�m�,~s����2���ܝMM
��,=?�d���&�t�{#	�x�}������ݼ��s�G���>�9��l�?3X�`���%]]��ToHA �I��)���W�w��fDv���k�#?
]w<�9w55^Ftw⪞mf��j�Txk^�a���~6�z�����ϲ��Vo[���˚����Z��m�����G�N�*J�X�$�@�J��L�jA��|�qG�U�I��O0Y�6j�"Hs�ĖYS⪞mf��aT��3G?�d���&�zY]�埅4`v�;w6s�O;,�	�@�	0[4>�3� �mKgՖ�K;e���"��u�֡�)�P<�N� �PmՂ��N ���i��vp��
4��`D�`�����DR���6a�*�(.�%HƔD:(�֥��ع��f�cT+��J�v�t��Ʊ�_�eD�Iїi��ݟ�^���\�}����}�8�YC�8����ۣ�P�Z]'\gWg��	�Z�kfc��2���8���+�^U�	Y���xjzӝ���I(͂��-����Zt%��m&<��dn��A�Z��m�YMdN�<@Iv��nt=:��:5A��p��$���͜P_�_S:g�RMm�o��'����Tj��^�G�E�BS�+��U�,�P!6���r����܌;���'����u��r��Zt%��m&<��dn��A�Z��m�YM|@յ�mDx�Ϝ��*@&��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M�"v�(=�@� �-k��R�	iT;��|B��2����&ՙ:Д;�d��nӸ{cDR���670��c%HƔD:(�֥��ع��������������Ʊ�_�eD�I�;��&��^���\�}]���!E�r &
�$J�� �X?�V޴�ik]�����4�;��|B��2����&�ۗ��/���د�гf[�?ez�@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�F�SZ�]b?,s�ca�s0CS� ��U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩ�JnFݲ��s����X�Q-�DAԄ��K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/8n
V~$�����1%��Ɇ�����5��Dao.\C�k]�	,��QUt�\��E;Eh	��V�>ȿ��'���#8=�<�^���pP�	ڹr����hi�aDU�G�a�E�}q^J=���ɛ�?өx(�i��/R�ݚ�Н�JnFݲ��s����X�Q�j*��{�%�@�V��l����,���R�e�0����[�4�f,o���
^���|6?������|�����X�Q����9gUS�|#9���
�:qEp�;�P�t�5fĉ>99��A0ok�׹��|�T��U�m7n,�
�$�P�����չ���1S������hi�aDU�G�a�E�נ���wf{��|6?���};4lW5�C�h\K�5~�o���sp%'�$x��9�&�P�w$��'HY-��Yk"1/o���sp%r�M$�*:���Z��b�8�dX��hWw�d�pP~��)%�����D��2E#fr�L�t�iZ]XF�hx��G��n����������������i�����d]���GF��a�1�Z���=�a�v��r��O}a �*/����k	�����}0x�'��D��ت��f��
i�c�r�h�5,Wlr�r%)cANU�:|��?�R��n���LH��BH�i	���P1�c8�Ŀ��s}��A��A�u�O}a 0=�.��4�� �����x?����Ji�];���IR*�fN�W�Ty��5�#�`���a��'�-
)\Y��?d��A �4<��!I�}Fh��K��dv��oTN֢&@��&̇i�d�?�-��i�m�T�੝�hy��Q�#<4^�H��bf�?ǉ�=�չ�Ad���&I���<�,���E�f�?ǉ�=ʘۥ<3�\�%�	V���W���Bm�����rk�[b�0<��-�����*���}�gf�mk�$���]׽��X;p`��D�����M�;��i_2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��"/���]�Q诤�e��C�`�/�t��cm�@�ᩖ%�!����5��fH�6J)�s���-�)��|���=f�}��U�����̾0���;���˔����vg�ĝ����a��X`��_/��;�y/Ә���@�ۻ|2���̂; ,@�� د<�l雲	k����ۥ�Y�m�չ���1�]����71d�G�E�y���(%��}kutC������i{�W�G��!?�d���&�C#/<���q��3�*�M}x�C���Q�$�SE��'HY-m�@8��/=�e���-��FG�n�t�iZ]XF�hx��G��!�`�(i3�(}y��������i�?d��A ��+���LQ�f�?ǉ�=G&%	��ڏ�<
DN��І��%n3������0�O���]�|��T�5�d�,W�hQ�GvE��?��%��h�r�|6�gb��A�h��+FeA'�u���}| �e����kn4@Q�/�!�`�(i3k/�z�xEQ���*[UxG!�`�(i3���ꀍ�˺�Q���f�?ǉ�=��9��稕C��S�w��iY�;����2��}��CϾH�)�h��=;�)�^�\q�\E��0ס�Wd�#jsrCm�k��/z*x�n;��|B_�&F���b?,s�ca�$G1�O�P�9�L�,���F@;��7,������Z�׽�刍X��!���ū���t�T��?E-h��`f���sC>��ӚH�RtV�^�'ž1�|�'����u��r��q�\E��0���ɥ�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r��pT/�GS�)���܇�a��o��ё\Bk�	�Ni�{�����f[*b~*��s��,l����M?��y�!�`�(i32W���R0(|v��t�a�^��D���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M|]η��q��_N�����,�ǰTm�v��G�g�v��Z�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U�Z�@ns䟳��LQ�%�+2��k��kK�I�Q4p�/Cj���C�1,�A��#�jV�{+��i�Iu�5�O�%E#P_TR�\+�[�ƪe�0cwU�R?�[6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3e�v��ҵl�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r��pT/�GS��%�����d��-��![L��^C�+a��o���H�RtV�^�3��C���H�� �YߥթD�[*�Bi�v�V��'�njVfV:)��{D~�u��r��!�`�(i3e�v��ҵl+��%�k<.�B�0���;�¬pX��g��U-�e�,���6+����%>�rGO�D mWN!�`�(i3�v�Wס���G�K$x/��&���Xd	�/I%L�Q��T��� h�ҩΪ���l�� m.x��(��p���'jsrCm�k�J��6�d�C�
���W��3��ݪ��=��l�r|{�,��5�Q�J��6�d�.�B�0���;�¬pX��u]9�#�I�s)l໶�,!�`�(i3�W�7�tM���p���'jsrCm�k�J��6�d�C�
���W��3��ݪ��=��l�r|{��\��~U�J��6�d�.�B�0���;�¬pX�出����mo�B� �b��!�`�(i3?V��j�c�:#��XB��4,�Q��U����z~��6��	���`y����ݚ�Н��Ra])n#���r����!�`�(i3:8�zH_ɗ�;2V-W��	c@�^ k�1{&��� M?��y�!�`�(i3!�`�(i3e�v��ҵl�]�!��	Ǹ�y85����[��xԲ ._�U6�bL�f�z�����jV�{+�fbmDF�!�`�(i3՝� s�#���k$ !�`�(i3{k�h�+&k@C�Ɨ0z�cULE��K3�j�U�V������:��`6;�¬pX���O��R�^Ƒ�ӆ�v�9��!�`�(i3��Ě�����}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j���_J��`U�a�(��^GѬ�_aT��3G?�d���&�����t���B8궩�t&%�=:���'��-�3��#?1�U���gFck
����ɣ�<�f��jV�{+��i�Iu�5�O�%E#P_TR�\+�[8$u�Ӵ-����t�T��?E-h��`f���sC>��ӚH�RtV�^�'ž1�|�'����u��r��q�\E��04>^!b!4b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3��Nh�=f[���������<�.�����8��GM��-����!�`�(i3e�v��ҵl�]�!��	Ǹ�y85��r��3��kO��u�+�uB;y�cU�^.����P�7� �:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6�8���SY�N�xʫ�A���;_��8W�w��fD)��J(�92�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�D� �B���9�V��r"nq���z���;�Ӏ�K��tV�:V%�&)�򄭩I4��欱���j�����|��ȤDL�>5�C����A��,��I4��欱���j�����s�QN���d���!it�td���52�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��Pdl2����}*X�K{�(��	}�@�r�<Uee�N�����0�=��;��|B���r�����z� 3P���@{2귑����Sa�!�`�(i3!�`�(i3���i����k]m����}Dq�f��z� 3P���@{2귑����|�kI��RhF��U>V%`�~�߇���t�k]m���E�i�m}66j�"Hs�@��C�,ԭ}3Y�Z��E��3?�d���&�Û=�������fo��ZpW4%"������k�I��RhF�䦓����������A2wKaC�IX0F�MV�ҁGG��Ւ��n�0 zK<U|r���3f�\�J��ײjw�ME�po守�ubs��2[�a��o���H�RtV�^����lr�{��|e��0�U+�qbp@���\ Nhk+Q�h'�Ȝx�5W ��̫(� h�ҩ���fCI��8��GM��-����<�6�Q=�I��� g~��q6g�yF}���V6l;�<��'�̗����Ep� �����4br���^��D�Ϛ�-����!�`�(i3�Y�
 �vc�jj&��G�9m6�̟�1��"~6���aq��3=]��m�D��-����!�`�(i3-3!E!����Bf���̓@?5ɔ��,Vr!�`�(i3��Id�!�`�(i3�XW�����5=��)Q���nF���<�W�.�P�	��
�Q�}<�6�Q=���F��O��ݚ�Н�烉s)�v�bP�63Z�t��Qѳ$G��A0ok��烉s)�v�T����� Ԕ׹�ն'�U;|�� �Rɮ�/���¨}�n/�J����lh�o��_�Rv�䩲$��ƣ�Ę�2{y����i�q,?5q�+�#4��F��8M�po守�ubs��2[�a��o���H�RtV�^��KV�9�]Kߩ�d��my$�N��o�/���;�I��Yq0�ʂ�j�Ï��	�l�lM�3 H�RtV�^���9���LQ�/81tSjv��� л��"�Nm>Ǖ��U�._�3
�v�v-}�	mp
���U{���8^��hJL��;���N�4��N	�7q������O�޳!?�R��n}�����H�X��WG ���N��b���c]p�5�	$o��Z�_�n�To�[�}�~��lg�7&�oe�XƤ5_���M���R��ӟ-���J��RQH�RtV�^�XW�����ZRR���dN�<@Iv��nt=:��:5A��p�I��Yq���k$ �� л��P�궊�2�����8!��?V�&�2���)x�?{���x.�Knq��5+*��4br������Ľ����Չxv��Օ��qvdЧ^{�j����'�����Z>ؼ��XyH�RtV�^<�6�Q=닓.�`�33c=��u<Rleށ�!�`�(i3��Qѳ$G��A0ok�®� л��5ߧE4��<�6�Q=���F��O�C#/<���q�5ߧE4���Qѳ$G�φ��<�6�닓.�`�3����΅�yǐ:�̋�:.�{��T����.������胋�M��a�-V�Cp	��?�?"���і�O:찹��S>���P��Y1C8�L�-�zm�2����~8GJ8���,�I}�F�y�^	#�-w˕���k�S���ld �jX��b�����ݻ��"~6���aq������J�?�d���&��������꓂O�q��.�1�4�o� c ��*�O.�N��A$�P������5d�������)G�9�=�1��*�
�I(͂X��WG ������&�Ko���&�@�}7�q��J��v1a{J�h�µj�!{�N<'��Il��!yZ�d/�����C�V���3��ֳ�Ե�i ӫ/��mR�MP��G�>��jj��r����.�aq���XF;�p)��
ۼ���Xv�"�M�)u��)o�0�ʂ�j�Ï��	�l�lM�3 �\Bk�	y�}�6f&r#o�]�ʄ�q������O�޳!?�R��n}�����H�X��WG ���?�,t�J�}D՛��W;���\�H��/Sg�w��'o�MdGN�������m��8\�Ia#i��N�Na����g�6���Q,|��,�ϣ퉧:��oQ�|i��N�Na����g�6���Q,|h���fn�g��]�J*�Rs�08�b(�����̜�I0���ԏ�.fOe	�HlU�!=���~�����gn�=4�4�	���WdM4@�肥�J����V��)x�?{���x.�KnqH�Ћ�r��%�z�J��z[�A���3�L����e�eV�M�z$��P�!�A˪[	��j"jȩ�i��N�Na����g�6���Q,|h���fn�g��]�J*�Rs�08�b(��R����� ӫ/��mt���������m���šB)��zR���b�3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$A�׭�%*b�3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�/%\��jX�m ޶&�hbvk~�#x�%��4�w����m�����F��O�n���šB)�X[��:~6q���w�=��u���'b�'=�(J�}�֖��-�X]t$IDW��E��q��u���'b�'=�(J�}�֖�
�c���zU���̜�I0���ԏ�.fOe	�HlU�!=���~�����gn�=4�4�	���WdM4@�肥�J�h@I �y ӫ/��mR�MP��GX��WG ���zR���b�3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�V�һ�d�#P�j2E�?��Id��o<Z�L5a�"Pn��s�I���I�����OeU���(;)(F�T��̙�R��I���I�����OeU���(h�a��Mg.6�k���'���o|k�Lb���'���o|k�Lb����k��?�,t�JN��	�Ȓ�cЉ�M�K���]��i�a�sir��5��܊K�+���w�PjI^�UI0���ԏ�.fOe	��<������r���3�:�����{~㽕���䕽v1a{J��=t�z/�����C�V���3�O��+�El�n�.��ɠ4�04�jf�nٚ�2�,�n�.��ɠ4�04�jfc¦�.��aY8.���׹��*P�{��	�ɭ��
/��y;��=�m�W��n4p�`6j�"Hs��Z�W����/��hH�C�F?�������L�����%C1��,2�A���ۖ��S�<Ԣ�,
�u#���n=�Z��W/��WuB=�r����'����IX0F�MV�ҁGG��ABk@�0h�5eצ'ž1�|�'����Ut�\��3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�V�һ�d�f��xp�M�C�x!�H�k��^)ҠN�2$�I))����A�m�(�}gQp�3+�\�G�����dc�@c�����hX��WG ���͹�k�9��d��-��!�L�F.	-�L��&PY~�y����o)�T*�c��܍w�S}�u��XC���}D՛��W;���\�H��/Sg�w��'o�MdGN����9�d�L�c]p�5�	$o��Z�_�n�To�[�}�~��l c�o�u��.ᬵy��o"#}aUt�\������-�G�h��\`�R�kA7��V ��݇!�
D���;�g��ޙVb�"�I���I�����OeU���(;�~1��_���̙�R��I���I�����OeU���(�&�r^-���.������v�8:������fI��jÇ+�_�n�To�[���9�P�4vE7�MW�o�>>����I���I�����OeU���(�G%i��A!��: ��ao.\C�kG��R�	J_g()��ikp���H���F��kt'n
V~$����4~V��3�L����e�eV�M�z$��P�!�A˪[	��j"jȩ�i��N�Na����g�6���Q,|h���fn��0h���J*�Rs�08�b(��un��7� ӫ/��mt������q�)]Q�x��r_��mzf	�$NT�I���I�����OeU���(;)(F�T��̙�R��I���I�����OeU���(h�a���4�M1��A���ۖ�k�V\�#P�j2E�?�5ߧE4��>je`��@d:�����{~�Vb�"�I���I�����OeU���(;)(F�T��̙�R��I���I�����OeU���(h�a��:��O�?�I))����A�m�(��C��AF�Р=��'e����&�@�}7�q��J��v1a{J�h�µj�!���5��Dao.\C�k]�	,��QUt�\�u��a��i��N�Na����g�6���Q,|��,�ϣ��19TH���"L?�����G�\�4���gn�=4�4�	���WdM4@�肥�J��eqm����gn�=4�4�	���WdM4@�肥�J�:�D5��h7�xȀ��D׏�����Mp�-a�D͢q��`�L�5ߧE4��; T�����8��GM�v�]��1VTҝD!u�Z����pG�p�P�m��������a-6�Da�K:+>N��	�Ȓ�cЉ�M�K���]�����` ��y/�����C�V���3��ֳ�Ե�i ӫ/��mR�MP��G���:��KY�[b%Ɨ����7�P�K�+���w���řA{���C�x!�H����'^_J���|{�mdJ�1���)�@����p�-a�D͢fU�9�׏�����MFi��|F�}�WP']��6�~����0D�N( Q���L}��M�~�ajJɫ �~wS �X�C���������C��֑xGV�eU���(;)(F�T�	�_��:��u���'b�'=�(J�}�֖�ت2�<�O��gn�=4�D-'��7�q����r� F�3N�����	��gn�=4�4�	���WdM4@��&����˶�ּX�b��c�fi�d\'�s�@#F e8�~����t9N\ا��=tu�㺅ڐK���l_��`N�z��7|^���~�@3�$��I)p�z!��U	�`�o��_�Rv�䩲$��8��I��.��|ȃ�A(�c���_G��Hb�wd�#<����Tk�-������c�����B)|DՃ���lf^�;��C+�G~���M��Nv�*~A�,��`������]kK�+���w� �s		��N���u��v1a{J�@<}��A@g()��ikp���H���4�:s� �q��]���~��-Y[;�wQ���սv1a{J��z*  x�I))����A�m�(���}܁'�O��<��J*�Rs�08�b(��l`��\1S�u{hK�'��݉�=�����w�=��u���'b�'=�(J�}�֖��-�X]t$I$�D���O�J*�Rs�08�b(��p�QD�á��&�@�}7�q��J��v1a{J�}D7B��#��M��hbD��ڙ�n�ZLN�	���}���x�A���ۖ��1�:��^ K=�b��ġ��,��{�	���v�8:?�'���&!����-�g()��ikp���H���G6.�~�݊���w�=�����C��֑xGV�eU���(;)(F�T�@Z
��#���Fi�"τ�����p��}��aq����(
}���û��i��N�N-��;��M�z$��PКą���g�U4���Z�Ϥ�h��K�r�\E�6O:��2bv!nU��K.��QW�4��i�P�
ɴ��z�4�	���WdM4@���d5���J*�Rs�08�b(��R����� ӫ/��m� ����+��J>�߯�"5�o٥眣TFC�)x�?{���x.�Knq��п��Tg()��ikp���H���G6.�~�݊��n����,6��œ�'�����Rkj}kq�MT�5�o[�a��[�s���J��sr�l�k]m��8����`�'J*�Rs�08�b(��R����� ӫ/��m� ����+��J>�߯�"5�o٥����Y�JM�b��v݋N�����7u7҃Q*�6������1�R+-h]�83NI�����w/,g{Y#0����l��=5; �e�W|��6�C��(3��7�q��J������-VL�Q�K��x�A���ۖ��S�<Ԣ�ɨ]^(���Ѹ���_�j�`���: ��ao.\C�k���uf|ò���
��_������B�K��1��n�da�ۣqM��X�~ ӫ/��m�D�K����g1�#�(�>^�l��e�eV�>�3�eZ~�f�R�&Aju�j[����#��47�
ɴ��z�D-'��7�q�����*8���������@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*�Va�ir�4br���qP�V>t'�̗����S]�_�_��Ut�\��"�Nm>�DQrv����)�x�.���;���8$_Z
��9�#���F�H۷`n
V~$ą�m[���'���c�e�+���4.�*�l��=5;�a���8n
V~$� ����%��>M���b��v݋N�����ה��#m��`$�\�����ZLN�	���nE�g%�zR���bJ�%Ph�r^m"�OB7A�SW�N����4�P��/ ں4��VJΣ8��3�L����e�eV�M�z$��P�!�A˪[	��*3)�����3�L����e�eV�M�z$��P�!�A˪[	�2��h�d�)x�?{���x.�Knq��!cI͸I))����A�m�(��C��AF�Р=��'e����&�@�}7�q��J��v1a{J�}D7B��#��T��n ^��A���ۖ"'��&އp��;�{����G�\�4���gn�=4�4�	���WdM4@��&����˶O@�s��M���c�v�J��sr�l�k]m��n���=�y���5Lwn�3
�v�v-}�	mp��"����I0���ԏ�.fOe	�HlU�!=T۳�͕��~K
eڟ7���&�@�}7�q��J��v1a{J�}D7B��#��.M�LYq^���&�@�}7�q��J��v1a{J�}D7B��#�w���{,�:g()��ikp���H���y���@�Krw�&�z<a�4�ڈt�[b%Ɨ���û��i��N�Na����g�6���Q,|]���#��:��oQ�|i��N�Na����g�6���Q,|6.o�7�OY����A�b��v݋N�����|�+��)�Р=��'e����&�@�}7�q��J��v1a{J�}D7B��#����5��Dao.\C�k]�	,��QUt�\�zf	�$NT�I���I�����OeU���(;�~1��_��pPo��zT۳�͕������4~V��3�L����e�eV�M�z$��PКą���gƜ*3)�����3�L����e�eV�M�z$��PКą���gơ��^��Mrw�&�z<a�4�ڈt׏�����MJ�1����z%�ژ�(�*4��%�#o�]�ʄ�q�����Q%I4��뇿D!�0�?�R��n}�����H�X��WG ��W|��6�C��(3��7�q��J������-VL�*3)����#�(�>^�l��e�eV��_�vԡ3�OY����Ag{Y#0����l��=5;N�����O������Mc�WT�D�3����K�F��_�M8O؏����:�~�1ߩ���ZAL�:������`4��D-~nҙ��ș5*�M��1�y�I��m�n����[�s���J��sr�l�k]m���������N��-���'�[�s���J��sr�l�k]m��M�s�Ӟ*��"xC��-�T(u	M^)FU9����8BW�R7���r_��m��zb����2�ę�u'b�'=�(��$��O
ɴ��z�4�	���WdM4@�p�r5A��J�1�����u���"6ɲ�cz���Ӵ�"�6j��;٬sf.���Y�m��
ɴ��z�4�	���WdM4@�݆M�g���󑟇���-hbvk~�#x}���y�Db��E(�\�H��/Sg�w��'o���u���"6����׾dC�ڃ�P �J�bMfo{��M�M������W&Z)�8�i{2!�Mn�g�L�2w�f��8/���u"MP�UUc�WT�D�3����K�F��^VE����t]���|���N(�1[�G���Kn��ɲ�cz���Ӵ�"�6j��;٬sf.���Y�m��
ɴ��z�D-'��7�q�������Q�$Gu�w��Ds��>���R�^J|WQ	��2�b��v݋N�����|�+��)�Р=��'e�C��(3���-��w��k]m��8Sg��
Ԧ�C��u����1m�Ut�\�8�%<}���"'��l������O05 S�s�lɲ�cz���ł)w���m�±��m|�b��Č�?��|��袔MUt��!�J��Y��̵�"xC��-�T(u	M^��|A�I���pP�$D\��z�
ɴ��z�4�	���WdM4@�E�RN�- \C��(3���-��w��k]m��������C��uu8I#M{c�}���Fo|k�Lbx(�i��/R�;b�-�2�׏�����M�[�S�n�H�,l�����(4G��>�S���%��V�c��ݕZ����pG�p�P�m�������3�� �f������.S��X��덎a-6�Da��J6����"'��l����C1zhi�Y
�,�LٗH�1�"'��l����C1zhZVv ?JZ��,H���F�]	
~ao.\C�k�Y�\�n����[�s���_����J������ݱ�JGy�ˆn����N��+�CAƨ�D5���a-6�Da��zb��B�>��֑xGV�05 S�s�l�1Qa����˓#�������\|u='�c�-��;��>�3�eZ~����z
��|u='�c�-��;��b'�Y@%^~>��mJ�1���K���L���4�04�jfx(�i��/R}�	76�&�� Ӗ�t$�)�vxv���}�_�� �R�"�n)�Q��ܾ7�'��ܷh������{ԕ����D#8`�k]m��v��z_����6��Ɔ ���Ve��˅�:�}��E5��OP�Յ������ꏶ�Ij�'��щĽ��1{�K�f(&�/� s�Y�����0�;�s�$�������E2��W䁱3�}$}��î�Zq�������L`G�v�~��]X���k���_��&7��N:��"^���H> �([�4����tm+�E^J*�Rs�08�b(������T���n��<��%m�Y$� 1���!��|�+4K-��4~H�<�&��x����<�S���c�&����:)x�?{���x.�Knq��5+*�����˱f�렾����o0hp�J$!@S�@��NXA��� �h��N�Mܲ���C�>5�,}9P!��|����GuDc%^oe�Y��k���_��&7��^�F��vh^���H> �s�bͦ-(�Ⱥ�kJ��*���[�\#���Ƹ��p��6�>������n�O��Ե�Z+���g��o����>�/�d�@���G3��X&+M?�n��<��%m�Y$� 1Z�����j�r]��=�찺pl�E(��6�� ~^N�gG`	Plh�P	���Mcyö��]f�,"y���L? ���U�d�@���GU����N�="��u���܁�i��:ژ�����Z4GL�}�痽�����)�aO��������J�)��Z+���g��o����>�/�d�@���G�%�4�'S!��#����В�S���GuDc%^oe�Y��k���_��&7��^�F��vh^���H> �ݎ' w%g��_���cشŀ��`�z���xl%����v缐%�/�<�|K7�&^v� E#�F2~��E,};�^�)׶9�H*.埲���G4��cf�l6�L� *���˿O�F�{�e4���ҏ�n�%$3��)�M8��	��?�'��/2RIh���o��G9�}Q*%΢Ӟe�H5��M���*�f;!+�+$�����^/e��d]� ���_�hbvk~�#x��q��ZVT�x�"��XƤ5_�J�	�LÆ���#��}���![<"XC}ץE�$��Ly����:�����U��2�ڥ����Ⱦ|����?��eߍ��鋎Z O\������U�._�nQ�rV��q�t7�.��/��SB�/���\VO�l� mr�m� Z�l�o����>�/�d�@���G�X���.��ġ��,l5R?}�b�+��z���&�2���)x�?{���x.�Knq���'
�?��p��6�>z8^�G8Lu�>�� 6�o8:4�I���c�90��c��qq:Fa�7���W"�P�K��q��[@��'ž1�|�'�������H��e��k�J��ֽ�\����g��U-�e>� {�}���my$�N���Uە��jz�\=�/��8y����Y)�'�m���[�4�f,�{_8�Y��=�}�Vݨ��\9�oA�d��JXl'�T��~��Uг�|<������M���LQ�/8n
V~$�+�$�i4�ǖ��`Y��}�O���硙�t�\������n�O��Ե�a(􆿳�e�&���6�+�$�i4�� N٣��}�O���硙�t�\��������J�)��a(􆿳�e�&���6�5ߧE4��J�1���k_���b_���~�L*f3�~�;kΗ�31���鸗r�!��=cv6�Ɛg)x�D�����X�X� U�X���#g�k����?��j:���'�Ȳ��A$�P������5d�B� ��~��U��B��-ն'�U;|=�9U'��A(�c���_G��Hb=��"�ԭ��\VO��1��0����,?}�a�,��Sq'�@8�Qq���z���nF���<�W�.�P��c3��4br�����w������n�5�����}�pIɽ�Jz_�b_X�XV�b�z'hۉ)K7͍���E@�����s��U;4���^a�nu4Bޗ��jw�	����/�ciJ��Yu�����Fodً]�N� &p�ۻ�F'i0QW��8�	3i�\��׹��t�M��|S�/���[�4�f,.�q����e8�b,Qk^|�ˮ���$:N�t%��zxa(􆿳�e�&���6A�іx���\&<���٘ۼ�%6Y�G�˱�ߓC娤l��
�~�qYUS���%��(ݒ�hU�y�搲)���$:N�t%��zxMg.6�k�5ߧE4��rw�&�z<a��N� φ��<�6��PT�!�wd�1�D�V��	��y����U����鸗r?1��j�=�*%΢Ӟe�a�f+(��R}��ک��\VO�l� mr�m�(�s׷�~O���M3X/��A���-�Vb� ���������J�)��a(􆿳������>�,r�/<]mz�(�����2a� `�ئ��# ��6U(�<"��q�
�`�N�9�;�S��2a� �6�_��f�D�!$9�:�A��� �c�eC(�5_��&7��Ј-�S��f~��DV��O8Ľ-�X]t$I��6U(�<"f6�8Nn.�!�6UVo��6U(�<";�~1��_�u�9j7Zj�� N٣���RUt�E��6U(�<"�; Me~��?���J��J�)����ʨ )o�or�K��:8���+����d�]�����0\)����+�ڔ�I�����t�a,�$a���h�4h;D8���:���`�����O�Y�a�G�'������E�n���
Ո�C�hk��Y��A�m�(�,"��h�2
��F�l��=5;z��˻N�dLd�r:ha3B��*w���6b��ʏ��Z��4`��O::��n[I?��8y����i��?}�˼�f���MWdWV��	��y��I�A���U2�h=c��_���	���%�� U2�h=c���9�Y��v�c��Q��"��0��C��-���R��)�xQ�b��v݋N������Q���u��N�"9���b�=�`~G��?.�#g�k��֓&Zf��%j_H�ˉ���0����f�Nd+l�Yҽ֗�x�\c�5#�y�mDƝ��0vdL�_E�������,�ǰ	M,��rER)�H[ɳv��X�x�LV(<���wj-�::��n[I?����$ڑ�N�(]n�5+�D�k�x<C��:�c-yi"�����2�^˧��t]����ض?l�� *%΢Ӟe�a�f+(����&�K�VF0��<�@QQO�W;D�gL4�e�d�Jw��3�	[ZZ��-�`��W��D5�|��7�OT�,���q5�n-�@�4ڧ�<�j�k�����Z���%�d��:
�r" ���]'\gWg��	�Z�kfc�L�C���e��S�J\7!c�2�����U��\ڦ'ž1�|�'����Ut�\��3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�nR��ړC娤l����pQ�q��!W�{_8�Y����X���������4~V��3�L����e�eV�M�z$��PЄ� *��eR��n�J>|�
#�`�^{��u�oDb_X�XV�b�z'hۉ)Ժ=���]��4br��L��_��R��n�J>|�
#�`�^{��u�oDb_X�XV�b�z'hۉ)K7͍���E@�����s��U;4���^a�nu4Bޗ��jw�	��#.w^�oG��8��GM/f��Z�~K
eڟ7���&�@�}7�q��J��v1a{J��(O T'Q`���$���^��y6�T���1���A%�@* ����c�v�J��sr�l�k]m��^~W���\'P�����M@�qX�Uu�T��3���W
�����4~V��3�L����e�eV�M�z$��PЄ� *��eR��n�J>|�
#�`�^{��u�oD�g�)�I�졉�&�@�}7�q��J��v1a{J�9�+J!��Q`���$���^��y6�T���1�����@�g����Ǵ=O�W;D�1X�iRd��D�����X���*"��Zʊӽ�����4br���v���R��n�J>|�
#�`�^{��u�oDE���7t�x(�i��/RŻ�&ǥ��a���F߸��S�Ȍ�w��ڷ�"�l�7%�]X����Ǵݵ��O��M`(繉�i�O��M`Օ���4���M���o�G�m�?���bq��;��|B���l
����>Ź9f���D5�|��7�OT�,	3i�\��׹��t�uDh/P^s[xkx U�_@�M��8S.�U��)���Y;e�iK ����)c���[�����3fEa�F��x�ޝE��A(�c���_G��Hb��a-6�Da�Ɔ ���/r�G�vH��~�.G�`��ٞ�R̕q������鷂�nF���W�_te*�"��?�.>#�����c�v�_����J����肥�Jӳ��n�5�����}�pIɽ�Jz_�b_X�XV�b�z'hۉ)Ժ=���]�X�C���������C��֑xGV�eU���(�˃��'�	3i�\��׹��t˔R��}K7͍���\C�
<r�8����H�v�ov�*�Y�G�˱�ߓC娤l��(Q6D���硙�t�\K7͍��|��W&":nv�q����� N٣�SG㴊�?����q5�n�JrPQV��dh_��tCdN�<@Iv��nt=:ྵp�!���k+Q�h'�Ȝx�5W ��̫(��a-6�Dae<�Ia��l�9W�a��=2oΠ�5�Y� u/2v:�v�H|���}�pIɽ�Jz_ꛨg��U-�eQ��,��ǖ��`Y�SG㴊�?����q5�n��dq�8���/�#P�j2E�?��6U(�<"e��w^9u�R̕q���s���4���܂%j_H�ˉE���Z�Y�G�˱�ߓC娤l��°������R�wX��)C8�o���C�x!�H��Tp�����5���7�~���=���q5�n�>.U$�o�N��	�Ȓ�cЉ�MMe9���ݱy�搲)���$:N�t%��zxMg.6�kzf	�$NT�I���I���C1zh�6���Q,|�b��暴�~���=���q5�n�>.U$�o��	�_��:�����C��֑xGV�eU���( �H^䁭	3i�\��׹��t�{ƨ��;N��-���'���c�v�_����J�����&����˶���n�5�����}�pIɽ�Jz_ꛀg�)�I�졉�&�@�}�-��w��k]m��n���=�y�y�搲)���$:N�t%��zxMg.6�kx(�i��/R#k�˟ܒ�o|k�Lb��ܐ�}�|&�xVgY��m������L}�E�6�����>Ź9f�Ps_*�GqW�w��fD`���$� �O"�2|�x�'�{��|�t3�e���S2�>��,+$\�M��ࣣ�{
��lҷgᗄ�xl��]���ҏ$ ~x==u�l��~	��c'PV�����[�'��#��ee[V	Q���7�5�h�5,Wluϛ�?udF���ˏ��Z���G�dE�h�����RyX�K{�(U4��\r�<Uee���R�}vJ^��u�*��?�d���&���}�7�v�k]m��7���
�Gbh��,������0��/������-Ӥ�v��د�r�QA�ј�;-;*�7�����G3҇
I��)���W�w��fD�Ɔ ���:U����w�R���y��E ��M�ee[V	Q��W< �mP�9ǧjK�|�� �2*�,��M���HaU$kX��@�?J`�p1��^���f��5��܊�W�-�4pm�|2;$�JأͽgF"?h�5,Wl�/�O'�=��#W�U���1��^���f��5��܊�iA'R�	�)l8�u0�P"G�wk����xC�(������Q�N��	�Ȓ��1��p3I��P`�k�)V��B�1/�����ٗ���3����,�ǰ��#x$E�ee[V	Q����de�ݤ��|�D+��V��m�̖˄��O�]�0=�f�U����*@mj�)�G�O\f��,+��(Pd��'�\#�5�'���I���y�c)�h�<om����4�&����Z�׍�R��ƿ;W ��.���:�Nz�]'\gWg��	�Z�kfc�_	�Ƽ���8|bs��2[�a��o���H�RtV�^�d�@���G�M��hb�Nҷ`=�}�Vݨ�W��]���uc��̄T�٥��TУ��xۛ�>�u��8�x�iH3�=���B���ꡝ���#RuZ��D�"����DZ�NU�=��1�������g�Z��3��a���!@�f")u��r��܌;���'����u��r��#�աl����aGl�97��EN�y�JB���PY~�y����o)�T*�c�Q��Ne<��t��7 �E�!6\|����?��������J*�Rs�08�b(����:����
�ݚ�Н���te�*EB�̟�1J�	�LÆ���#����-/a8!�`�(i3���8�2����o�W��g��Ȋ�>�������Ra])n#���r������{$@d�̟�1���	���#!�`�(i3�5ߧE4��9�d�L��d�@���G-*��j�J�	�LÆ���#����-/a8!�`�(i3���8�2N5�Hɫ'���+m�ol��Ә�~1S�vw�b!�`�(i3��jVѭ@!�`�(i3��i��}�12�mj�{�N<'��I!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍu���q�_/;W ��.���)�2�r;��|BL˓ }4o�X�G[��l÷{H�D�d�@���G��3v�qnQ�rVY���K*�O���t�h���rg���̟�1�w�H�-4b��he=��$M��J���]�Yl;��|B�A�ω�K��� �R�QبM��u!/��"�*�����M���R��ӟ-���4�&����Z��hs������No�ߏ�����"?��A$�P������5d�������y�(����<m�r$ɓǃl[�Ƶ�1tSjv��ߎ ��E�5���u�L���nF���<�W�.�P��c3��4br��yO{��`�
n��>�my$�N��]流�>���ݤ�E��p�����-i�q ���$5�nc�Gy=��g����Ǵ=q@L����F��� ��f�{_8�Y��=�}�VݨuN�wAB��O���&z�вԺL�9�T�I����y���c��ᥟB�'��a�S���%�����ռt
�AԢ�a\蟟Q��ǺΕR��ӟ-�q�x�~<��w���	�e�<j��.#՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r��;�jmT�#�YN
��)e���^b�~H����8�O�5���1tSjv�!�`�(i3�YN
��)e������p�r~�h��ݚ�Н���w�w:�!�`�(i3%Q�[�J����˦G�K7͍��|��W&":�ݚ�Н�$f��_Ub�F�S�1 ��H�����4br��>�=,W�[�?�R��n}�����Hٚ�-����!�`�(i3	�)��&ghRV��R�4br���h�Һ�!�`�(i3��jVѭ@!�`�(i3	�)��&ghRV��RK7͍��|��W&":�ݚ�Н�$f��_Ub���r�������W��{��I�+��X��WG ��hw�U�1S���%��V�c���Ǵc�1�RG�p�P�m��������a-6�DaA�іx�~=&lL�i ����yw�kkr��;���};#P�j2E�?��˓#����j�V܎L��dE��İ���K7͍��|��W&":�xȀ��D׏�����Mp�-a�D͢q��`�L�x�$�M���)���߄�	�\M?��y���L�ΪA��YN
��)e�*8Җ�N��k�=H����8�O�5���n
V~$�j�V܎L������ⰷ���4br��$��x�-O��T���B�R���>_��\��;}{�t���=�gdN�<@Iv��nt=:�z�X
3kZ�x(�i��/R�P�HS|�O�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�k��{`.~��No�ߏ��T�4(���;��|BJ�U�� �X�G[�wE�=p���4br����3v�qh�5,Wlr�r%)cAQ17�b�����d���!i�/��mS%rƂ�o��+rp�叧���5ʦ���'�QV[1��<[��a�D��<F��� ��f�{_8�Y��=�}�Vݨh��J)7�������<�02r��dN�<@Iv��nt=:���/z*x�n;��|Bʦ?�H#F`�� �R�ćTm���j��u�Nb#¯��TG6�o8:4�I���c�90��G��6�(&�L��'ž1�|�'����u��r�������i҆�w��kf�6�(�A?'���c�e�|E��΢�Mr��p�ԍ�S��4$:��{K·��ΥT�tE�ŀ�sb�*� �XU�*��l�lG�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G����l�� U�9��n	-�L��&PY~�y����o)�T*�c���&����ŷ�k��d䖬n���S滑����ZLN�	���:����
�K:+>�͵�p۱e��0���J*�Rs�08�b(��MdGN���!�`�(i3�a;���a��Bf���͵�p����#�=3!�`�(i3��˓#��͚��m�Bx&����˦G�����"�fĉ>99��A0ok��fĉ>99��o|k�Lb�"������U�._�h�5,Wlr�r%)cAH�Ћ�r�H�RtV�^�G:w��-6�$�Dr��c<.~\�H��/Sg�w��'o�MdGN���!�`�(i3
x�ߜ�BɆJӱ�zW,D#kZ_�U2����}Dq�f��	��x���"n�Κ�-6�$�Da��Q����ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�Sm�6��`4�04�jf�*4��%�#o�]�ʄ�	�)�N�O�W;D�0gv�%Z?�R��n}�����H�-M�O��~��rpf�2&tRW��n
}vh�xC��f0� �-:���h��e�z����,_�k������I�3���o��(fw���'�̗������O�j�v�Ut�\�� ����%��>M����?"3�m�����h�n*��(� �C� �1�����Ǹ���)/�~�T���]�q9+t�}8BW�R7���r_��m>f��8�D�u��u���)������x�ԉ�>x(�i��/R&����1㋾����IdN�^�%��>M��_L�"����A|�stUy��{oFU�b�$��Ut�\�� ����%��>M��_L�"����A|�stUy��{o@�f�WfTUt�\�2b���J����w_���!�b[�Mv!���xB�R���>_��.�2��0tNF5��q���v�{n��뾦�c�}���Fo|k�Lbx(�i��/R�;b�-�2�׏�����M�[�S�n�H�,l����M?��y��W)�x�F[�-6�$�DK�(+�`W��,8���|b�,�ۮAH�œ%�	�)�N�	-�L��&PY~�y����o)�T*�c�p��;�{��,"�~�K���9��4�Ä/�,o� �ҋ�;��.�[ ٓ���p��e�_y.O�%T��C�~0ޭ�A|�stUy��DbY}n��!g�θ�8���d�W�J��H����8�(����X��WG ���4O/3�L�3B�\G��C.mg��n��뾦�p�-a�D͢q��`�L�N�]�B���vE���GFOg�S�<�c�!���X���z�`�|e�3B�\GJ�8;��w�h��Jc'�yK�w���"X��[��Q[R�7HN��R��bP�63Z�t�5ߧE4��Fr��jCZ�zk��X���#7�I�Jw��3�HU6�0�\��S��4$��}���`�|e�3B�\GJ�8;��w�h��Jc'�yK�w��
��Q�# 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��Wv�A����w�V�"~�ӵ(r7�8� ��$d������`7�tȈ������9P�-�,�AG�<���X饿��!�iv�aQ�Ϧ�M�ኾ���L��r�U���f��/?L���u�D��D1��n������� �k,
"i�̄�ѭ���ɿ�kF��l�l"��l䋬5Kq!�`�(i3!�`�(i3}��[b:��'(K�lc���97PC�e>2Tg�չ���1Y]H]w�
��P��*|��P�˩eNUD60L����q�?T���T��� ��?c�ĭႿ��h�q��r����$l�
�H�t���� *ί�$�E�#s�ss�7\�	�������;"��*G�e[u�;0�쒕��l\�����=@��Ù��\�����;��c���X��3i�+� a⣃_B�M�˵·�ۥ�Y�m�չ���1�]����7��j���N66j�"HsplS'yJ�p��)�}� ���x®�{9�%��t���8����Z��zH��\NیL_��f�Ä/�,o썀���P�e[u�;0��?w����3�s�'��U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩ�JnFݲ��s�5�>U�m�j*��{�%L_��f�����,���R�e�0����[�4�f,�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r���s�Yls��8��GM��-����!�`�(i3����]dF!�O+�|/������Lx�A�B��8�nb �z�g��U-�ew���7VaN�\�]
��s�G��38����]dF!�O+�|�����˨g��U-�e�,���6+�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ��R_�����xZ;a{-�X���!1B�0�/N�\�]
��s�G��38����]dF!�O+�|�ι�l�-䤔���8@[�_zβrE��g�Hbw���1����*����OE�)�%E��'Z*)�?�R��n��h
:h����t�h��W+��W��*#�m z����Z��oE�g�������(ӈ�����$��LSm�f�e8�1ޞ��&e[u�;0�2����k���RN�-#���$�m�7Y'��k���=R��Ԗ�A$�P������5d�C#/<���q{y����i�q,?5q��7���9��e���W� �{Z+ճpo守�ubs��2[�a��o���H�RtV�^�<��	B�ɔ9Q<ϯ)P<�ܓ�Y�� л�����g�Z��3��a���!@�f")u��r��;�E����=�O�-v�*_�mS8<�n�ݚ�Н�@20߀�����P0����3��x�p��!�`�(i3��&.��8�F�S�1 �烉s)�v�bP�63Z�t�u��I�Ɨy�"c�|����"�`��P��*|C#/<���qL��M����4�	��������A$�P������5d�C#/<���q{y����i�q,?5q�+�#4��F��8M�� л��'ž1�|�'����u��r���G��^���J��sr�lE�g�������(ӈ���m�r����I��Yq0�ʂ�j�Ï��	�l�lM�3 H�RtV�^R���Xc��Yu�����a��� vc�jj&��G�9m6�XƤ5_���"~6���aq���s{�'!�u��r��<�6�Q=2VP��Ѣ��P@JɈ.���3R��6 y2��R�\ Nh�;�P�t�5�� л��5ߧE4�흔\ Nh$�)�vx'X���5����'G�+p�9���?�(�JZ�Vk�;��|B��loXBȱg�S>X;Z�˯��R����e���Wƍ ٻ�l���M���R��ӟ-���4�&����Z��W�\7�(�ɔ9Q<ϯ���쨷	
P���ɒ�!�6UVo��`�m�;����^F�=�_�7V�o��_�Rv�䩲$����tb���~�26��\� :����JHn��z��r9�3C>��Ӛ��S�J\7CZ�zk��X��z�1P�үle�0��|#HK��A(�c���_G��Hb� h�ҩ�pi�NWHC�ۥ�Y�m/��kOT�����y������	SN��r�J��p��b���Nq#5z�dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3�#}�{��~v� 1��&k@C�Ɨ0z�cULE��K3�jAԢ�a\��ĂB/�缍kv޶Gla��Mp��֙l@�B�!�`�(i3�kv޶Gl���lr�q��p��b��������/!�`�(i3t�td���5;�jmT�#ʬw�S���d��-��!��EJ��7ޅ7�=w�'�̗����S]�_�_��u��r��!�`�(i3Sm�f�e�=�⳿P��}Dq�f���.J7h��,?��&�)�
�k\�i��}Dq�f��߆�p�h��{$�������LQ�/8۶&��L�H�W�J��H����8�O�5���1tSjv�!�`�(i3�Н��Ei1.��2����|e"�B�'��a���� Ev��\��;�,
�:qEp'{w#/ B!�`�(i3Sm�f�e8�1ޞ��&e[u�;0�2����k��d����j��8�u��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��}�6�nq�Z�@���v0��L�r:�}�6�nq�4�	��������A$�P������5d�C#/<���q{y����i�q,?5q�+�#4��F��8M�� л��'ž1�|�'����u��r���G��^���J��sr�lE�g�������(ӈ���m�r����I��Yq0�ʂ�j�Ï��	�l�lM�3 H�RtV�^R���Xc��Yu�����a��� vc�jjM�ｂ g�����j��8!��?V0D�	�I���_
�u�Y���H�hbvk~�#x�DS�AvF̓@?5�#j�o���&�2��������j���L�F.0D�	�I���_
�u�����|�G�p�P�C������H8Џ�Ӿ���yi�1tSjv����y��lD(�D �6�|�;�ƇT��J��sr�l�ԝy'��� л��5ߧE4��<�6�Q=���F��O�C#/<���q��ܐ�}ī:f����p��'G�+p�9���?�����,�ǰ����adp��e���Wƭ(n6eF�/�B|0<2��'7�u
f�.�c�n��`�7�,��n6�o8:4�I���c�90��G��6�iI9�o«IX0F�M�H{���<�e��BFbs��2[�a��o���H�RtV�^+���G����$�\%e��}Dq�f�#� �,W���Ǉ�y!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^i��H�p¢	�B�d���%������4s����ڕ3��t�ƍd��U>�Q�c6��?��!�6ʬw�S����}Dq�f��5ߧE4��"T^r��~����k�_�mS8<�nZ�~�|}�"����Ż�&ǥ��bP�63Z�t�5ߧE4��Fr��j��k���;V�
pFV�$=+R�˩��*��� ��U�_:�E��t?����a렾����޴8"��J�a$�Y �t/�(�P�KZ	��\#�Z¥���5.'MtZ�R����DZ��}�1U��VP\@Ww6CE!H^��Ƨ�0/��U��|:��'!�P�P2����+�wձ}���8y�����e�Q�� �)ԴG<�鶰.����܍ \O~��z����
����7,������Z�ך�>1Y�>c��?�B�t�xr�t��b����J�"I �����w���'�(�]�[�H���,&ǚ���φ��<�6�@a� ��fFMqlg��z?F�#��S�J\7O.�x�����(���2$�m�����G�'ž1�|�'����u��r��RD�~���M��V!�D��nF���<�W�.�P�	��
�Q�}g��A�L��d��JXl'�T��~��Uг�|<m�����G܌;���'����u��r�����Fz���2�b=���i�Wg�l���鯻��U��O�D mWNs_ѧ�p�O�D mWN���J�a��IX0F�Mb�Xϋ?@�n���/l�̬���	p|�O�E/�9��"J j�E��'Z*)�?�R��nj��P_Q����t�h��W+��W����uR���_�#g� |cz�����]X����7�4��~n�2o� �2�L2��R�͢��n-΂��m9Ϲ��*��x��� ���JH����8��#I�ND�s���H�V��-���^S��$�Gy��e���W������)<��U��)���Y;e�iK!���d."�9ŭ,iI9�o«IX0F�M��ŊPTWo9���b��|2;�E����A(�c���_G��Hb� h�ҩ�� ͷ�	���6�
V����b+}y[<�6�Q=�B -�6���'�QDndN�<@Iv��nt=:��:5A��p,�u�S��d��JXl'�T��~��Uг�|<!�`�(i3���9���LQ�/81tSjv����y��lD�TaDe��"�/֖�Yk{:fh�3�:5A��p�� л���������Z¥���5.'MtZ�R�!�`�(i3��&.��8�F�S�1 �烉s)�v�bP�63Z�t�u��I����~�Lk݁ 1���tw�i�Ք�w��y����J�a��?�d���&�J2���n�7�ct�����?
Z+6/Ahr����B�z���b�~8GJ8��"'���xO��H{��4-�9���{��Psmi'l:}��Q\�>�7���o��_�Rv�䩲$��V���,�wO0 zK<U|r���3fX�?���'��>��ԑ�%;�E����A(�c���_G��Hb� h�ҩ�h�x��JyW$q(W���ƍ2���l��^{T~H���^a�nu4Bޗ��jw�	���ݚ�Н���fCI��8��GMZ���Ӗ���mFA�$�!�`�(i3����,Ů�뒒���97��EN�fԯA&b닓.�`�3u���# �%��,�V�B�
X��Z����b�Ի�!�`�(i3�(��p�m���
y������Ľ���ANʂ'�8���y}	�'C�R7 �E�!6\
��7t��i��E�y�H�RtV�^߇�\���*���H��w�u�M�Һ����1)uם�!�`�(i3��&.��8�F�S�1 �烉s)�v�bP�63Z�t�u��I�Ɨy�"c���? 6����,�ǰx͝�I��D�X�����t<�NA��qޠ	S�uimK�ֶ����6�o8:4�I���c�90��6:����+�^n=\f�5>�I!�[�������QQ��B�"}��r$ɓǃl[�Ƶ�1tSjv���R�?�Γ�]#�y�W�CbE�{_8�Y��=�}�Vݨ��}Dq�f�S�#p���zՠ�����˦G�K7͍��|��W&":C#/<���q����g�Z��3��a���!@�f")u��r��R���Xc��Yu�������&G���y��lD���j��z$��
�5L��m}I������jH�2�s��� H���Y�����&G!�`�(i3�r���Ipˏ-).^QQBպW � ����i9v�I��`j!�`�(i3��&.��8�F�S�1 ��po守�uQw�$��Z��/�dW���3����V$=�b�oj�+p�K�J�iN�Sˇ^�6�H����8��� I���\�b��v݋N�����i�!w���p��;�{��!�`�(i3�<��	B��D厺��+�̟�14�����{��O?��ʔ��,Vr<�6�Q=��jVѭ@!�`�(i3S�#p���zՠ�����˦G�K7͍��|��W&":�ݚ�Н�烉s)�v�bP�63Z�t��Qѳ$G��A0ok��烉s)�v�T����� Ԕ׹�Ӫ��*$���A�<M��[��k�}�t��/�dW�<龈��ơlП���V03Y��9�`�I��W����Ľ��M�ȅõ����(�x�HM���#g�s�
�`�I��W�^��D����jVѭ@���Fz�!�`�(i3!�`�(i3S`�@�4:��]�����n�h��N�M��~��f�!���zՠ�~��q6g�yF}���V6l;�<��'�̗����#!d�+I0���ԏ�.fOe	�N:w�h?Y�)�}���"���d����yi�l,V�,k� sȸ�"rR!�`�(i3�����z�>9G`�(���'�5�,�xs�*"1���)�=�w�������:�5}`'l:}��Qb!��u����$A�O1�Et�]�!����M[��Ǣs��j�ŉ��m�n�~�!�G���-7s�9���o>��l%i�-�F*D@��j�i�p��+��~���O!��Q]� _ό���.��|�����E ����7dh�?зq8�Ј'���Xw�,bxqX�b!��u�<�`A��_i3i 
�c��]�!����M[��Ǣs��j�ŉ�|�w��DK����$���7s�9���o>��l%i�-�F*D@��j�i�p��+�/s�1��p��Q]� _�rs�i���`�M�	=̞��>��3
�v�v-}�	mp,��_А#�<om��F`���G���`y���C#/<���q�5����`KiW��
�!C� �u؅��FJ��gm?2�I��6�]���~`��ʿ��^�����èV�H�?���E�m ��?Z��G.�w�v�d����x�l��1:�N�*�x�� л���D��������m#p�W��	]�	M$E�Z�ݚ�Н����iYM�5q{! l��2
L./;�Ly�Af�?ǉ�=񔿄�aB6Э~���V��2
L.�X;p`��3
�v�v-}�	mp,��_А#�<om���'$W$�X�<�6�Q=�L�K��%<7�`+Al��R��������,NL ���<�6�Q=�o�f�Ԝe���b�!�`�(i3�(�;\��B�}�ݚ�Н��D���R]���gRI/!�`�(i3X&|a�#g()��ikp���H������7Pr��ġ��,�&�C�/�s�f�I��b��v�#$�q�
k-���w�E�V{�!�`�(i3�V�����/>�"�Ax!�`�(i3��3�N;C�]�'!�`�(i3�7Z.m�w��'�k�f!�`�(i3�u~xgA���������6%�a�k���n�}�� �с�'(�U�c�&8�,��
�Q!}-[BvGޣkQ�A���ۖ$����nQ�rV,?�����ݚ�Н��43S�d��ރ;�{��C�{����K�7��C4%̈́��� л�6�R�W� W��|E�q��w\F�M$E�Z�ݚ�Н�H���!�>�*�!�`�(i3���K�7��8C+a�Rj�~���0ȓM�Me��^��>�z'�:�N�*�x�� л� ��$�,���X;p`����$AA�:JϮ����j���ӱ}�tM�@;w�$C,0�?���<�6�Q=4?s����k-����b=�<�6�Q=�0V32;5�-�����4)cq�vG+|�<�� л����ٜ�]�X;p`���C�,�4���y��lD�Vf�`H�j��-@��ey�E���x�ր�ݚ�Н��y�3���k�K��hczZ����4b�zvѓ�!�`�(i3�7?�S�!!�`�(i3�$�~c/~�O��������y��lD�Vf�`H�jT��b9���ey�E�����$���f�?ǉ�=A#�
�v!�`�(i3��%ў׫=�F�K�@�!�`�(i3V��uL$��!�`�(i3�$�~c/v��&EA)�� л�֕ߝԀ�#kcBTX�#�
�ge[I��4�	����������P�=��:F�|���m�:�-22�v ,��rQd->�d�!�`�(i3f�������9�|Nb��'1-�,bxqX��ƿ�d���5�[՚1D��c�e��o����B��7dh�?��,:&���z2%警�d��]�Q��f�_��BvGޣkQ�A���ۖ$����nQ�rV�}!�@�?0d׻zc��7U�	Y���۠ql��*O��_^=�/Jt\�J���70�'���O�V2y/�ߓ��y��]��K��Xw�e60�' ��[w�{0
����)��#L����?;����IX0F�MV�ҁGG`5:��0}}��*ꅺS�J\7�p���"Z�v��!<�6�Q=�r$ɓǃl[�Ƶ�1tSjv��� л��	�%1A��b+}y[��\ Nhk+Q�h'�Ȝx�5W ��̫(� h�ҩγpo守�u��"����G��Hb� h�ҩή� л��	�%1A�qo<�khku��J�>�V����f�z��SR:g()��ikp���H������7Pr��ġ��,�i�/Q�ಧ�y��lD&[�x�R�"��}Dq�f���&.��8�}Q�sd��]� )�+��p���"��NwK�"&'��Y_�C#/<���qH^��Ƨ�0	�Ʊ�R���uoJ`AP�n�M�t䖬n���S滑����ZLN�	���<~=��<��?6Ґ�6�d45sf��ݚ�Н�<�6�Q=��b+}y[R��X鷴QW�w��fD!J��/٣׆p�9��+:��0	��